-- generated with romgen by MikeJ
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity CG_BASIC is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of CG_BASIC is


  type ROM_ARRAY is array(0 to 16383) of std_logic_vector(7 downto 0);
  constant ROM : ROM_ARRAY := (
    x"F3",x"AF",x"C3",x"74",x"06",x"C3",x"00",x"40", -- 0x0000
    x"C3",x"00",x"40",x"E1",x"E9",x"C3",x"00",x"00", -- 0x0008
    x"C3",x"03",x"40",x"C5",x"06",x"01",x"18",x"2E", -- 0x0010
    x"C3",x"06",x"40",x"C5",x"06",x"02",x"18",x"26", -- 0x0018
    x"C3",x"09",x"40",x"C5",x"06",x"04",x"18",x"1E", -- 0x0020
    x"C3",x"0C",x"40",x"11",x"15",x"40",x"18",x"E3", -- 0x0028
    x"C3",x"0F",x"40",x"11",x"1D",x"40",x"18",x"E3", -- 0x0030
    x"C3",x"12",x"40",x"11",x"25",x"40",x"18",x"DB", -- 0x0038
    x"C3",x"D9",x"05",x"C9",x"00",x"00",x"C3",x"C2", -- 0x0040
    x"03",x"CD",x"2B",x"00",x"B7",x"C0",x"18",x"F9", -- 0x0048
    x"0D",x"0D",x"1F",x"1F",x"01",x"01",x"5B",x"1B", -- 0x0050
    x"0A",x"1A",x"08",x"18",x"09",x"19",x"20",x"20", -- 0x0058
    x"0B",x"78",x"B1",x"20",x"FB",x"C9",x"01",x"18", -- 0x0060
    x"1A",x"C3",x"CA",x"05",x"31",x"F8",x"41",x"11", -- 0x0068
    x"80",x"40",x"21",x"F7",x"18",x"01",x"27",x"00", -- 0x0070
    x"C3",x"40",x"01",x"21",x"01",x"58",x"3A",x"80", -- 0x0078
    x"F8",x"CB",x"4F",x"20",x"09",x"22",x"A4",x"40", -- 0x0080
    x"CD",x"46",x"38",x"22",x"A4",x"40",x"21",x"E5", -- 0x0088
    x"41",x"36",x"3A",x"23",x"70",x"23",x"36",x"2C", -- 0x0090
    x"23",x"22",x"A7",x"40",x"11",x"3B",x"01",x"06", -- 0x0098
    x"1C",x"21",x"52",x"41",x"36",x"C3",x"23",x"73", -- 0x00A0
    x"23",x"72",x"23",x"10",x"F7",x"06",x"15",x"36", -- 0x00A8
    x"C9",x"23",x"23",x"23",x"10",x"F9",x"2A",x"A4", -- 0x00B0
    x"40",x"2B",x"70",x"CD",x"70",x"38",x"CD",x"8F", -- 0x00B8
    x"1B",x"CD",x"AF",x"06",x"CD",x"C9",x"01",x"21", -- 0x00C0
    x"18",x"01",x"CD",x"A7",x"28",x"CD",x"B3",x"1B", -- 0x00C8
    x"38",x"F5",x"D7",x"B7",x"20",x"13",x"21",x"00", -- 0x00D0
    x"40",x"23",x"7C",x"B5",x"28",x"1C",x"7E",x"47", -- 0x00D8
    x"2F",x"77",x"BE",x"70",x"28",x"F3",x"25",x"18", -- 0x00E0
    x"11",x"CD",x"5A",x"1E",x"B7",x"C2",x"97",x"19", -- 0x00E8
    x"EB",x"2B",x"3E",x"8F",x"46",x"77",x"BE",x"70", -- 0x00F0
    x"20",x"CD",x"2B",x"11",x"14",x"44",x"DF",x"DA", -- 0x00F8
    x"7A",x"19",x"11",x"CE",x"FF",x"22",x"B1",x"40", -- 0x0100
    x"19",x"22",x"A0",x"40",x"CD",x"4D",x"1B",x"21", -- 0x0108
    x"21",x"01",x"CD",x"A7",x"28",x"C3",x"19",x"1A", -- 0x0110
    x"4D",x"45",x"4D",x"20",x"53",x"49",x"5A",x"45", -- 0x0118
    x"00",x"43",x"4F",x"4C",x"4F",x"55",x"52",x"20", -- 0x0120
    x"42",x"41",x"53",x"49",x"43",x"0D",x"00",x"FF", -- 0x0128
    x"FF",x"FF",x"C3",x"6B",x"01",x"C3",x"4F",x"01", -- 0x0130
    x"C3",x"5D",x"01",x"1E",x"2C",x"C3",x"A2",x"19", -- 0x0138
    x"ED",x"B0",x"21",x"01",x"C0",x"3A",x"00",x"C0", -- 0x0140
    x"B7",x"C2",x"7B",x"00",x"C3",x"8B",x"00",x"CD", -- 0x0148
    x"83",x"01",x"3E",x"01",x"07",x"10",x"FD",x"0F", -- 0x0150
    x"47",x"1A",x"B0",x"12",x"C9",x"CD",x"83",x"01", -- 0x0158
    x"3E",x"FE",x"07",x"10",x"FD",x"0F",x"47",x"1A", -- 0x0160
    x"A0",x"12",x"C9",x"D7",x"CF",x"28",x"CD",x"83", -- 0x0168
    x"01",x"E5",x"1A",x"1F",x"10",x"FD",x"21",x"FF", -- 0x0170
    x"FF",x"38",x"01",x"23",x"CD",x"9A",x"0A",x"E1", -- 0x0178
    x"CF",x"29",x"C9",x"CD",x"1C",x"2B",x"FE",x"08", -- 0x0180
    x"D2",x"4A",x"1E",x"F5",x"CF",x"2C",x"CD",x"02", -- 0x0188
    x"2B",x"F1",x"47",x"04",x"C9",x"FF",x"FF",x"FF", -- 0x0190
    x"FF",x"FF",x"FF",x"FF",x"FF",x"D7",x"E5",x"3A", -- 0x0198
    x"99",x"40",x"B7",x"20",x"06",x"CD",x"58",x"03", -- 0x01A0
    x"B7",x"28",x"11",x"F5",x"AF",x"32",x"99",x"40", -- 0x01A8
    x"3C",x"CD",x"57",x"28",x"F1",x"2A",x"D4",x"40", -- 0x01B0
    x"77",x"C3",x"84",x"28",x"21",x"28",x"19",x"22", -- 0x01B8
    x"21",x"41",x"3E",x"03",x"32",x"AF",x"40",x"E1", -- 0x01C0
    x"C9",x"3E",x"1C",x"CD",x"3A",x"03",x"3E",x"1F", -- 0x01C8
    x"C3",x"3A",x"03",x"ED",x"5F",x"32",x"AB",x"40", -- 0x01D0
    x"C9",x"3A",x"1C",x"43",x"EE",x"01",x"D3",x"FF", -- 0x01D8
    x"32",x"1C",x"43",x"C9",x"3A",x"27",x"44",x"EE", -- 0x01E0
    x"0A",x"32",x"27",x"44",x"C9",x"D9",x"06",x"08", -- 0x01E8
    x"16",x"00",x"CD",x"FA",x"01",x"10",x"FB",x"7A", -- 0x01F0
    x"D9",x"C9",x"C5",x"DB",x"FF",x"E6",x"01",x"5F", -- 0x01F8
    x"DB",x"FF",x"E6",x"01",x"AB",x"1F",x"30",x"F8", -- 0x0200
    x"3C",x"AB",x"5F",x"3A",x"12",x"43",x"47",x"10", -- 0x0208
    x"FE",x"DB",x"FF",x"E6",x"01",x"AB",x"CB",x"22", -- 0x0210
    x"B2",x"57",x"C1",x"C9",x"CD",x"1F",x"02",x"D9", -- 0x0218
    x"F5",x"0E",x"08",x"57",x"CD",x"D9",x"01",x"3A", -- 0x0220
    x"10",x"43",x"47",x"10",x"FE",x"7A",x"07",x"57", -- 0x0228
    x"DC",x"D9",x"01",x"3A",x"11",x"43",x"47",x"10", -- 0x0230
    x"FE",x"0D",x"20",x"E8",x"F1",x"D9",x"C9",x"06", -- 0x0238
    x"FF",x"3E",x"AA",x"CD",x"1F",x"02",x"10",x"FB", -- 0x0240
    x"3E",x"66",x"18",x"D3",x"E5",x"D5",x"C5",x"21", -- 0x0248
    x"69",x"35",x"11",x"00",x"00",x"3A",x"23",x"40", -- 0x0250
    x"5F",x"19",x"7E",x"32",x"26",x"F0",x"32",x"27", -- 0x0258
    x"F0",x"01",x"AA",x"80",x"CD",x"FA",x"01",x"B9", -- 0x0260
    x"20",x"F7",x"3E",x"FF",x"A9",x"4F",x"10",x"F4", -- 0x0268
    x"CD",x"FA",x"01",x"FE",x"66",x"20",x"F9",x"3E", -- 0x0270
    x"2A",x"32",x"26",x"44",x"32",x"27",x"44",x"C1", -- 0x0278
    x"D1",x"E1",x"C9",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0280
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0288
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0290
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x0298
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x02A0
    x"FF",x"FF",x"FF",x"FF",x"CD",x"14",x"03",x"22", -- 0x02A8
    x"DF",x"40",x"CD",x"E2",x"41",x"31",x"88",x"42", -- 0x02B0
    x"CD",x"FE",x"20",x"3E",x"2A",x"CD",x"2A",x"03", -- 0x02B8
    x"CD",x"B3",x"1B",x"DA",x"66",x"00",x"D7",x"CA", -- 0x02C0
    x"97",x"19",x"FE",x"2F",x"28",x"4F",x"CD",x"4C", -- 0x02C8
    x"02",x"CD",x"ED",x"01",x"FE",x"55",x"20",x"F9", -- 0x02D0
    x"06",x"06",x"7E",x"B7",x"28",x"09",x"CD",x"ED", -- 0x02D8
    x"01",x"BE",x"20",x"ED",x"23",x"10",x"F3",x"CD", -- 0x02E0
    x"E4",x"01",x"CD",x"ED",x"01",x"FE",x"78",x"28", -- 0x02E8
    x"BB",x"FE",x"3C",x"20",x"F5",x"CD",x"ED",x"01", -- 0x02F0
    x"47",x"CD",x"14",x"03",x"85",x"4F",x"CD",x"ED", -- 0x02F8
    x"01",x"77",x"23",x"81",x"4F",x"10",x"F7",x"CD", -- 0x0300
    x"ED",x"01",x"B9",x"28",x"DA",x"3E",x"43",x"32", -- 0x0308
    x"26",x"44",x"18",x"D6",x"CD",x"ED",x"01",x"6F", -- 0x0310
    x"CD",x"ED",x"01",x"67",x"C9",x"EB",x"2A",x"DF", -- 0x0318
    x"40",x"EB",x"D7",x"C4",x"5A",x"1E",x"20",x"8A", -- 0x0320
    x"EB",x"E9",x"C5",x"4F",x"CD",x"C1",x"41",x"3A", -- 0x0328
    x"9C",x"40",x"B7",x"79",x"C1",x"C3",x"64",x"05", -- 0x0330
    x"FF",x"FF",x"D9",x"F5",x"CD",x"33",x"00",x"CD", -- 0x0338
    x"48",x"03",x"32",x"A6",x"40",x"F1",x"D9",x"C9", -- 0x0340
    x"E5",x"2A",x"20",x"40",x"11",x"00",x"44",x"B7", -- 0x0348
    x"C3",x"D9",x"04",x"FF",x"FF",x"C3",x"9D",x"30", -- 0x0350
    x"CD",x"C4",x"41",x"D5",x"CD",x"2B",x"00",x"D1", -- 0x0358
    x"C9",x"AF",x"32",x"99",x"40",x"32",x"A6",x"40", -- 0x0360
    x"CD",x"AF",x"41",x"C5",x"2A",x"A7",x"40",x"06", -- 0x0368
    x"F0",x"CD",x"D9",x"05",x"F5",x"48",x"06",x"00", -- 0x0370
    x"09",x"36",x"00",x"2A",x"A7",x"40",x"F1",x"C1", -- 0x0378
    x"2B",x"D8",x"AF",x"C9",x"CD",x"58",x"03",x"B7", -- 0x0380
    x"C0",x"18",x"F9",x"AF",x"32",x"9C",x"40",x"3A", -- 0x0388
    x"9B",x"40",x"B7",x"C8",x"3E",x"0D",x"D5",x"CD", -- 0x0390
    x"9C",x"03",x"D1",x"C9",x"F5",x"D5",x"C5",x"4F", -- 0x0398
    x"1E",x"00",x"FE",x"0C",x"28",x"10",x"FE",x"0A", -- 0x03A0
    x"20",x"03",x"3E",x"0D",x"4F",x"FE",x"0D",x"28", -- 0x03A8
    x"05",x"3A",x"9B",x"40",x"3C",x"5F",x"7B",x"32", -- 0x03B0
    x"9B",x"40",x"79",x"CD",x"3B",x"00",x"C1",x"D1", -- 0x03B8
    x"F1",x"C9",x"E5",x"DD",x"E5",x"D5",x"DD",x"E1", -- 0x03C0
    x"D5",x"21",x"DD",x"03",x"E5",x"4F",x"1A",x"A0", -- 0x03C8
    x"B8",x"C2",x"33",x"40",x"FE",x"02",x"DD",x"6E", -- 0x03D0
    x"01",x"DD",x"66",x"02",x"E9",x"D1",x"DD",x"E1", -- 0x03D8
    x"E1",x"C1",x"C9",x"CD",x"AF",x"06",x"3A",x"80", -- 0x03E0
    x"F8",x"FE",x"12",x"20",x"0D",x"CD",x"A9",x"38", -- 0x03E8
    x"3A",x"40",x"F8",x"CB",x"57",x"28",x"F9",x"CD", -- 0x03F0
    x"B0",x"38",x"21",x"36",x"40",x"01",x"01",x"F8", -- 0x03F8
    x"16",x"00",x"0A",x"5F",x"AE",x"73",x"A3",x"20", -- 0x0400
    x"10",x"14",x"2C",x"CB",x"01",x"30",x"F3",x"3A", -- 0x0408
    x"80",x"F8",x"CB",x"5F",x"C2",x"D4",x"04",x"AF", -- 0x0410
    x"C9",x"5F",x"21",x"18",x"40",x"3A",x"80",x"F8", -- 0x0418
    x"CB",x"4F",x"C2",x"C9",x"04",x"CB",x"67",x"C2", -- 0x0420
    x"D0",x"04",x"3E",x"07",x"BA",x"28",x"E8",x"7A", -- 0x0428
    x"07",x"07",x"07",x"57",x"0E",x"01",x"79",x"A3", -- 0x0430
    x"20",x"05",x"14",x"CB",x"01",x"18",x"F7",x"3A", -- 0x0438
    x"80",x"F8",x"47",x"7A",x"C6",x"40",x"FE",x"60", -- 0x0440
    x"30",x"13",x"CB",x"08",x"30",x"31",x"C6",x"20", -- 0x0448
    x"57",x"3A",x"40",x"F8",x"E6",x"10",x"7A",x"28", -- 0x0450
    x"26",x"D6",x"60",x"18",x"22",x"D6",x"70",x"30", -- 0x0458
    x"10",x"C6",x"40",x"FE",x"3C",x"38",x"02",x"EE", -- 0x0460
    x"10",x"CB",x"08",x"30",x"12",x"EE",x"10",x"18", -- 0x0468
    x"0E",x"07",x"CB",x"08",x"30",x"01",x"3C",x"21", -- 0x0470
    x"50",x"00",x"5F",x"16",x"00",x"19",x"7E",x"21", -- 0x0478
    x"18",x"40",x"CB",x"76",x"28",x"24",x"FE",x"2B", -- 0x0480
    x"38",x"20",x"FE",x"30",x"30",x"04",x"D6",x"2B", -- 0x0488
    x"18",x"16",x"FE",x"3B",x"38",x"14",x"FE",x"5B", -- 0x0490
    x"30",x"04",x"D6",x"36",x"18",x"0A",x"FE",x"60", -- 0x0498
    x"38",x"08",x"FE",x"7B",x"30",x"04",x"D6",x"3B", -- 0x04A0
    x"C6",x"C0",x"32",x"24",x"40",x"57",x"01",x"00", -- 0x04A8
    x"20",x"CD",x"60",x"00",x"7A",x"FE",x"0D",x"28", -- 0x04B0
    x"07",x"FE",x"01",x"28",x"03",x"C0",x"EF",x"C9", -- 0x04B8
    x"21",x"18",x"40",x"CB",x"B6",x"FE",x"01",x"18", -- 0x04C0
    x"F4",x"3E",x"40",x"AE",x"77",x"AF",x"18",x"DD", -- 0x04C8
    x"CB",x"FE",x"18",x"F9",x"3A",x"24",x"40",x"18", -- 0x04D0
    x"A6",x"ED",x"52",x"11",x"28",x"00",x"B7",x"ED", -- 0x04D8
    x"52",x"30",x"FB",x"19",x"7D",x"E1",x"C9",x"79", -- 0x04E0
    x"B7",x"28",x"3E",x"FE",x"0B",x"28",x"0A",x"FE", -- 0x04E8
    x"0C",x"20",x"1B",x"AF",x"DD",x"B6",x"03",x"28", -- 0x04F0
    x"15",x"DD",x"7E",x"03",x"DD",x"96",x"04",x"47", -- 0x04F8
    x"CD",x"29",x"05",x"20",x"FB",x"0E",x"0A",x"CD", -- 0x0500
    x"3C",x"05",x"10",x"F4",x"18",x"16",x"CD",x"29", -- 0x0508
    x"05",x"20",x"FB",x"CD",x"3C",x"05",x"FE",x"0D", -- 0x0510
    x"C0",x"DD",x"34",x"04",x"DD",x"7E",x"04",x"DD", -- 0x0518
    x"BE",x"03",x"79",x"C0",x"DD",x"36",x"04",x"00", -- 0x0520
    x"C9",x"3E",x"07",x"D3",x"F8",x"3E",x"7F",x"D3", -- 0x0528
    x"F9",x"3E",x"0F",x"D3",x"F8",x"DB",x"F9",x"E6", -- 0x0530
    x"EF",x"FE",x"2F",x"C9",x"3E",x"07",x"D3",x"F8", -- 0x0538
    x"3E",x"7F",x"D3",x"F9",x"3E",x"0E",x"D3",x"F8", -- 0x0540
    x"79",x"D3",x"F9",x"3E",x"07",x"D3",x"F8",x"3E", -- 0x0548
    x"FF",x"D3",x"F9",x"3E",x"0F",x"D3",x"F8",x"AF", -- 0x0550
    x"D3",x"F9",x"3E",x"0F",x"D3",x"F8",x"3E",x"01", -- 0x0558
    x"D3",x"F9",x"79",x"C9",x"FA",x"1F",x"02",x"C2", -- 0x0560
    x"9C",x"03",x"C3",x"3A",x"03",x"31",x"F8",x"41", -- 0x0568
    x"AF",x"D3",x"FF",x"21",x"00",x"F4",x"11",x"01", -- 0x0570
    x"F4",x"01",x"FF",x"03",x"36",x"00",x"ED",x"B0", -- 0x0578
    x"0E",x"FF",x"ED",x"78",x"E6",x"08",x"47",x"D3", -- 0x0580
    x"FC",x"ED",x"78",x"E6",x"08",x"21",x"11",x"37", -- 0x0588
    x"11",x"00",x"38",x"A8",x"00",x"00",x"D3",x"FD", -- 0x0590
    x"ED",x"78",x"E6",x"08",x"21",x"69",x"35",x"A8", -- 0x0598
    x"18",x"12",x"D3",x"FE",x"ED",x"78",x"E6",x"08", -- 0x05A0
    x"21",x"0A",x"37",x"A8",x"20",x"06",x"21",x"31", -- 0x05A8
    x"37",x"11",x"23",x"38",x"E5",x"EB",x"11",x"F0", -- 0x05B0
    x"42",x"01",x"23",x"00",x"ED",x"B0",x"E1",x"11", -- 0x05B8
    x"90",x"43",x"01",x"10",x"00",x"ED",x"B0",x"C3", -- 0x05C0
    x"6C",x"00",x"AF",x"D3",x"ED",x"3A",x"04",x"F8", -- 0x05C8
    x"CB",x"57",x"C2",x"00",x"00",x"C3",x"C0",x"06", -- 0x05D0
    x"FF",x"E5",x"3E",x"0E",x"CD",x"33",x"00",x"48", -- 0x05D8
    x"C3",x"00",x"30",x"FE",x"20",x"30",x"25",x"FE", -- 0x05E0
    x"0D",x"CA",x"62",x"06",x"FE",x"1F",x"28",x"29", -- 0x05E8
    x"FE",x"01",x"28",x"6D",x"11",x"E0",x"05",x"D5", -- 0x05F0
    x"FE",x"08",x"28",x"34",x"FE",x"18",x"28",x"2B", -- 0x05F8
    x"FE",x"09",x"28",x"42",x"FE",x"19",x"28",x"39", -- 0x0600
    x"FE",x"0A",x"C0",x"D1",x"77",x"78",x"B7",x"28", -- 0x0608
    x"CF",x"7E",x"23",x"CD",x"33",x"00",x"05",x"18", -- 0x0610
    x"C7",x"CD",x"C9",x"01",x"41",x"E1",x"E5",x"C3", -- 0x0618
    x"E0",x"05",x"CD",x"30",x"06",x"2B",x"7E",x"23", -- 0x0620
    x"FE",x"0A",x"C8",x"78",x"B9",x"20",x"F3",x"C9", -- 0x0628
    x"78",x"B9",x"C8",x"2B",x"7E",x"FE",x"0A",x"23", -- 0x0630
    x"C8",x"2B",x"3E",x"08",x"CD",x"33",x"00",x"04", -- 0x0638
    x"C9",x"3E",x"17",x"C3",x"33",x"00",x"CD",x"48", -- 0x0640
    x"03",x"E6",x"07",x"2F",x"3C",x"C6",x"08",x"5F", -- 0x0648
    x"78",x"B7",x"C8",x"3E",x"20",x"77",x"23",x"D5", -- 0x0650
    x"CD",x"33",x"00",x"D1",x"05",x"1D",x"C8",x"18", -- 0x0658
    x"EF",x"37",x"F5",x"3E",x"0D",x"77",x"CD",x"33", -- 0x0660
    x"00",x"3E",x"0F",x"CD",x"33",x"00",x"79",x"90", -- 0x0668
    x"47",x"F1",x"E1",x"C9",x"3E",x"08",x"D3",x"FF", -- 0x0670
    x"32",x"1C",x"43",x"21",x"D2",x"06",x"11",x"00", -- 0x0678
    x"40",x"01",x"36",x"00",x"ED",x"B0",x"3D",x"3D", -- 0x0680
    x"20",x"F1",x"06",x"27",x"12",x"13",x"10",x"FC", -- 0x0688
    x"21",x"AB",x"34",x"11",x"50",x"43",x"01",x"38", -- 0x0690
    x"00",x"ED",x"B0",x"3E",x"01",x"32",x"14",x"43", -- 0x0698
    x"21",x"30",x"39",x"22",x"8C",x"43",x"21",x"DB", -- 0x06A0
    x"39",x"22",x"8E",x"43",x"C3",x"6D",x"05",x"3A", -- 0x06A8
    x"00",x"C0",x"FE",x"43",x"CA",x"01",x"C0",x"3A", -- 0x06B0
    x"00",x"C0",x"FE",x"44",x"CA",x"01",x"C0",x"C9", -- 0x06B8
    x"3A",x"00",x"C0",x"FE",x"43",x"CA",x"01",x"C0", -- 0x06C0
    x"C3",x"AE",x"19",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x06C8
    x"FF",x"FF",x"C3",x"96",x"1C",x"C3",x"78",x"1D", -- 0x06D0
    x"C3",x"90",x"1C",x"C3",x"D9",x"25",x"C9",x"00", -- 0x06D8
    x"00",x"C9",x"00",x"00",x"FB",x"C9",x"00",x"01", -- 0x06E0
    x"E3",x"03",x"00",x"07",x"40",x"20",x"49",x"07", -- 0x06E8
    x"E4",x"30",x"00",x"44",x"01",x"01",x"03",x"06", -- 0x06F0
    x"E7",x"04",x"43",x"00",x"00",x"50",x"52",x"C3", -- 0x06F8
    x"00",x"50",x"C7",x"00",x"00",x"3E",x"00",x"C9", -- 0x0700
    x"21",x"80",x"13",x"CD",x"C2",x"09",x"18",x"06", -- 0x0708
    x"CD",x"C2",x"09",x"CD",x"82",x"09",x"78",x"B7", -- 0x0710
    x"C8",x"3A",x"24",x"41",x"B7",x"CA",x"B4",x"09", -- 0x0718
    x"90",x"30",x"0C",x"2F",x"3C",x"EB",x"CD",x"A4", -- 0x0720
    x"09",x"EB",x"CD",x"B4",x"09",x"C1",x"D1",x"FE", -- 0x0728
    x"19",x"D0",x"F5",x"CD",x"DF",x"09",x"67",x"F1", -- 0x0730
    x"CD",x"D7",x"07",x"B4",x"21",x"21",x"41",x"F2", -- 0x0738
    x"54",x"07",x"CD",x"B7",x"07",x"D2",x"96",x"07", -- 0x0740
    x"23",x"34",x"CA",x"B2",x"07",x"2E",x"01",x"CD", -- 0x0748
    x"EB",x"07",x"18",x"42",x"AF",x"90",x"47",x"7E", -- 0x0750
    x"9B",x"5F",x"23",x"7E",x"9A",x"57",x"23",x"7E", -- 0x0758
    x"99",x"4F",x"DC",x"C3",x"07",x"68",x"63",x"AF", -- 0x0760
    x"47",x"79",x"B7",x"20",x"18",x"4A",x"54",x"65", -- 0x0768
    x"6F",x"78",x"D6",x"08",x"FE",x"E0",x"20",x"F0", -- 0x0770
    x"AF",x"32",x"24",x"41",x"C9",x"05",x"29",x"7A", -- 0x0778
    x"17",x"57",x"79",x"8F",x"4F",x"F2",x"7D",x"07", -- 0x0780
    x"78",x"5C",x"45",x"B7",x"28",x"08",x"21",x"24", -- 0x0788
    x"41",x"86",x"77",x"30",x"E3",x"C8",x"78",x"21", -- 0x0790
    x"24",x"41",x"B7",x"FC",x"A8",x"07",x"46",x"23", -- 0x0798
    x"7E",x"E6",x"80",x"A9",x"4F",x"C3",x"B4",x"09", -- 0x07A0
    x"1C",x"C0",x"14",x"C0",x"0C",x"C0",x"0E",x"80", -- 0x07A8
    x"34",x"C0",x"1E",x"0A",x"C3",x"A2",x"19",x"7E", -- 0x07B0
    x"83",x"5F",x"23",x"7E",x"8A",x"57",x"23",x"7E", -- 0x07B8
    x"89",x"4F",x"C9",x"21",x"25",x"41",x"7E",x"2F", -- 0x07C0
    x"77",x"AF",x"6F",x"90",x"47",x"7D",x"9B",x"5F", -- 0x07C8
    x"7D",x"9A",x"57",x"7D",x"99",x"4F",x"C9",x"06", -- 0x07D0
    x"00",x"D6",x"08",x"38",x"07",x"43",x"5A",x"51", -- 0x07D8
    x"0E",x"00",x"18",x"F5",x"C6",x"09",x"6F",x"AF", -- 0x07E0
    x"2D",x"C8",x"79",x"1F",x"4F",x"7A",x"1F",x"57", -- 0x07E8
    x"7B",x"1F",x"5F",x"78",x"1F",x"47",x"18",x"EF", -- 0x07F0
    x"00",x"00",x"00",x"81",x"03",x"AA",x"56",x"19", -- 0x07F8
    x"80",x"F1",x"22",x"76",x"80",x"45",x"AA",x"38", -- 0x0800
    x"82",x"CD",x"55",x"09",x"B7",x"EA",x"4A",x"1E", -- 0x0808
    x"21",x"24",x"41",x"7E",x"01",x"35",x"80",x"11", -- 0x0810
    x"F3",x"04",x"90",x"F5",x"70",x"D5",x"C5",x"CD", -- 0x0818
    x"16",x"07",x"C1",x"D1",x"04",x"CD",x"A2",x"08", -- 0x0820
    x"21",x"F8",x"07",x"CD",x"10",x"07",x"21",x"FC", -- 0x0828
    x"07",x"CD",x"9A",x"14",x"01",x"80",x"80",x"11", -- 0x0830
    x"00",x"00",x"CD",x"16",x"07",x"F1",x"CD",x"89", -- 0x0838
    x"0F",x"01",x"31",x"80",x"11",x"18",x"72",x"CD", -- 0x0840
    x"55",x"09",x"C8",x"2E",x"00",x"CD",x"14",x"09", -- 0x0848
    x"79",x"32",x"4F",x"41",x"EB",x"22",x"50",x"41", -- 0x0850
    x"01",x"00",x"00",x"50",x"58",x"21",x"65",x"07", -- 0x0858
    x"E5",x"21",x"69",x"08",x"E5",x"E5",x"21",x"21", -- 0x0860
    x"41",x"7E",x"23",x"B7",x"28",x"24",x"E5",x"2E", -- 0x0868
    x"08",x"1F",x"67",x"79",x"30",x"0B",x"E5",x"2A", -- 0x0870
    x"50",x"41",x"19",x"EB",x"E1",x"3A",x"4F",x"41", -- 0x0878
    x"89",x"1F",x"4F",x"7A",x"1F",x"57",x"7B",x"1F", -- 0x0880
    x"5F",x"78",x"1F",x"47",x"2D",x"7C",x"20",x"E1", -- 0x0888
    x"E1",x"C9",x"43",x"5A",x"51",x"4F",x"C9",x"CD", -- 0x0890
    x"A4",x"09",x"21",x"D8",x"0D",x"CD",x"B1",x"09", -- 0x0898
    x"C1",x"D1",x"CD",x"55",x"09",x"CA",x"9A",x"19", -- 0x08A0
    x"2E",x"FF",x"CD",x"14",x"09",x"34",x"34",x"2B", -- 0x08A8
    x"7E",x"32",x"89",x"40",x"2B",x"7E",x"32",x"85", -- 0x08B0
    x"40",x"2B",x"7E",x"32",x"81",x"40",x"41",x"EB", -- 0x08B8
    x"AF",x"4F",x"57",x"5F",x"32",x"8C",x"40",x"E5", -- 0x08C0
    x"C5",x"7D",x"CD",x"80",x"40",x"DE",x"00",x"3F", -- 0x08C8
    x"30",x"07",x"32",x"8C",x"40",x"F1",x"F1",x"37", -- 0x08D0
    x"D2",x"C1",x"E1",x"79",x"3C",x"3D",x"1F",x"FA", -- 0x08D8
    x"97",x"07",x"17",x"7B",x"17",x"5F",x"7A",x"17", -- 0x08E0
    x"57",x"79",x"17",x"4F",x"29",x"78",x"17",x"47", -- 0x08E8
    x"3A",x"8C",x"40",x"17",x"32",x"8C",x"40",x"79", -- 0x08F0
    x"B2",x"B3",x"20",x"CB",x"E5",x"21",x"24",x"41", -- 0x08F8
    x"35",x"E1",x"20",x"C3",x"C3",x"B2",x"07",x"3E", -- 0x0900
    x"FF",x"2E",x"AF",x"21",x"2D",x"41",x"4E",x"23", -- 0x0908
    x"AE",x"47",x"2E",x"00",x"78",x"B7",x"28",x"1F", -- 0x0910
    x"7D",x"21",x"24",x"41",x"AE",x"80",x"47",x"1F", -- 0x0918
    x"A8",x"78",x"F2",x"36",x"09",x"C6",x"80",x"77", -- 0x0920
    x"CA",x"90",x"08",x"CD",x"DF",x"09",x"77",x"2B", -- 0x0928
    x"C9",x"CD",x"55",x"09",x"2F",x"E1",x"B7",x"E1", -- 0x0930
    x"F2",x"78",x"07",x"C3",x"B2",x"07",x"CD",x"BF", -- 0x0938
    x"09",x"78",x"B7",x"C8",x"C6",x"02",x"DA",x"B2", -- 0x0940
    x"07",x"47",x"CD",x"16",x"07",x"21",x"24",x"41", -- 0x0948
    x"34",x"C0",x"C3",x"B2",x"07",x"3A",x"24",x"41", -- 0x0950
    x"B7",x"C8",x"3A",x"23",x"41",x"FE",x"2F",x"17", -- 0x0958
    x"9F",x"C0",x"3C",x"C9",x"06",x"88",x"11",x"00", -- 0x0960
    x"00",x"21",x"24",x"41",x"4F",x"70",x"06",x"00", -- 0x0968
    x"23",x"36",x"80",x"17",x"C3",x"62",x"07",x"CD", -- 0x0970
    x"94",x"09",x"F0",x"E7",x"FA",x"5B",x"0C",x"CA", -- 0x0978
    x"F6",x"0A",x"21",x"23",x"41",x"7E",x"EE",x"80", -- 0x0980
    x"77",x"C9",x"CD",x"94",x"09",x"6F",x"17",x"9F", -- 0x0988
    x"67",x"C3",x"9A",x"0A",x"E7",x"CA",x"F6",x"0A", -- 0x0990
    x"F2",x"55",x"09",x"2A",x"21",x"41",x"7C",x"B5", -- 0x0998
    x"C8",x"7C",x"18",x"BB",x"EB",x"2A",x"21",x"41", -- 0x09A0
    x"E3",x"E5",x"2A",x"23",x"41",x"E3",x"E5",x"EB", -- 0x09A8
    x"C9",x"CD",x"C2",x"09",x"EB",x"22",x"21",x"41", -- 0x09B0
    x"60",x"69",x"22",x"23",x"41",x"EB",x"C9",x"21", -- 0x09B8
    x"21",x"41",x"5E",x"23",x"56",x"23",x"4E",x"23", -- 0x09C0
    x"46",x"23",x"C9",x"11",x"21",x"41",x"06",x"04", -- 0x09C8
    x"18",x"05",x"EB",x"3A",x"AF",x"40",x"47",x"1A", -- 0x09D0
    x"77",x"13",x"23",x"05",x"20",x"F9",x"C9",x"21", -- 0x09D8
    x"23",x"41",x"7E",x"07",x"37",x"1F",x"77",x"3F", -- 0x09E0
    x"1F",x"23",x"23",x"77",x"79",x"07",x"37",x"1F", -- 0x09E8
    x"4F",x"1F",x"AE",x"C9",x"21",x"27",x"41",x"11", -- 0x09F0
    x"D2",x"09",x"18",x"06",x"21",x"27",x"41",x"11", -- 0x09F8
    x"D3",x"09",x"D5",x"11",x"21",x"41",x"E7",x"D8", -- 0x0A00
    x"11",x"1D",x"41",x"C9",x"78",x"B7",x"CA",x"55", -- 0x0A08
    x"09",x"21",x"5E",x"09",x"E5",x"CD",x"55",x"09", -- 0x0A10
    x"79",x"C8",x"21",x"23",x"41",x"AE",x"79",x"F8", -- 0x0A18
    x"CD",x"26",x"0A",x"1F",x"A9",x"C9",x"23",x"78", -- 0x0A20
    x"BE",x"C0",x"2B",x"79",x"BE",x"C0",x"2B",x"7A", -- 0x0A28
    x"BE",x"C0",x"2B",x"7B",x"96",x"C0",x"E1",x"E1", -- 0x0A30
    x"C9",x"7A",x"AC",x"7C",x"FA",x"5F",x"09",x"BA", -- 0x0A38
    x"C2",x"60",x"09",x"7D",x"93",x"C2",x"60",x"09", -- 0x0A40
    x"C9",x"21",x"27",x"41",x"CD",x"D3",x"09",x"11", -- 0x0A48
    x"2E",x"41",x"1A",x"B7",x"CA",x"55",x"09",x"21", -- 0x0A50
    x"5E",x"09",x"E5",x"CD",x"55",x"09",x"1B",x"1A", -- 0x0A58
    x"4F",x"C8",x"21",x"23",x"41",x"AE",x"79",x"F8", -- 0x0A60
    x"13",x"23",x"06",x"08",x"1A",x"96",x"C2",x"23", -- 0x0A68
    x"0A",x"1B",x"2B",x"05",x"20",x"F6",x"C1",x"C9", -- 0x0A70
    x"CD",x"4F",x"0A",x"C2",x"5E",x"09",x"C9",x"E7", -- 0x0A78
    x"2A",x"21",x"41",x"F8",x"CA",x"F6",x"0A",x"D4", -- 0x0A80
    x"B9",x"0A",x"21",x"B2",x"07",x"E5",x"3A",x"24", -- 0x0A88
    x"41",x"FE",x"90",x"30",x"0E",x"CD",x"FB",x"0A", -- 0x0A90
    x"EB",x"D1",x"22",x"21",x"41",x"3E",x"02",x"32", -- 0x0A98
    x"AF",x"40",x"C9",x"01",x"80",x"90",x"11",x"00", -- 0x0AA0
    x"00",x"CD",x"0C",x"0A",x"C0",x"61",x"6A",x"18", -- 0x0AA8
    x"E8",x"E7",x"E0",x"FA",x"CC",x"0A",x"CA",x"F6", -- 0x0AB0
    x"0A",x"CD",x"BF",x"09",x"CD",x"EF",x"0A",x"78", -- 0x0AB8
    x"B7",x"C8",x"CD",x"DF",x"09",x"21",x"20",x"41", -- 0x0AC0
    x"46",x"C3",x"96",x"07",x"2A",x"21",x"41",x"CD", -- 0x0AC8
    x"EF",x"0A",x"7C",x"55",x"1E",x"00",x"06",x"90", -- 0x0AD0
    x"C3",x"69",x"09",x"E7",x"D0",x"CA",x"F6",x"0A", -- 0x0AD8
    x"FC",x"CC",x"0A",x"21",x"00",x"00",x"22",x"1D", -- 0x0AE0
    x"41",x"22",x"1F",x"41",x"3E",x"08",x"01",x"3E", -- 0x0AE8
    x"04",x"C3",x"9F",x"0A",x"E7",x"C8",x"1E",x"18", -- 0x0AF0
    x"C3",x"A2",x"19",x"47",x"4F",x"57",x"5F",x"B7", -- 0x0AF8
    x"C8",x"E5",x"CD",x"BF",x"09",x"CD",x"DF",x"09", -- 0x0B00
    x"AE",x"67",x"FC",x"1F",x"0B",x"3E",x"98",x"90", -- 0x0B08
    x"CD",x"D7",x"07",x"7C",x"17",x"DC",x"A8",x"07", -- 0x0B10
    x"06",x"00",x"DC",x"C3",x"07",x"E1",x"C9",x"1B", -- 0x0B18
    x"7A",x"A3",x"3C",x"C0",x"0B",x"C9",x"E7",x"F8", -- 0x0B20
    x"CD",x"55",x"09",x"F2",x"37",x"0B",x"CD",x"82", -- 0x0B28
    x"09",x"CD",x"37",x"0B",x"C3",x"7B",x"09",x"E7", -- 0x0B30
    x"F8",x"30",x"1E",x"28",x"B9",x"CD",x"8E",x"0A", -- 0x0B38
    x"21",x"24",x"41",x"7E",x"FE",x"98",x"3A",x"21", -- 0x0B40
    x"41",x"D0",x"7E",x"CD",x"FB",x"0A",x"36",x"98", -- 0x0B48
    x"7B",x"F5",x"79",x"17",x"CD",x"62",x"07",x"F1", -- 0x0B50
    x"C9",x"21",x"24",x"41",x"7E",x"FE",x"90",x"DA", -- 0x0B58
    x"7F",x"0A",x"20",x"14",x"4F",x"2B",x"7E",x"EE", -- 0x0B60
    x"80",x"06",x"06",x"2B",x"B6",x"05",x"20",x"FB", -- 0x0B68
    x"B7",x"21",x"00",x"80",x"CA",x"9A",x"0A",x"79", -- 0x0B70
    x"FE",x"B8",x"D0",x"F5",x"CD",x"BF",x"09",x"CD", -- 0x0B78
    x"DF",x"09",x"AE",x"2B",x"36",x"B8",x"F5",x"FC", -- 0x0B80
    x"A0",x"0B",x"21",x"23",x"41",x"3E",x"B8",x"90", -- 0x0B88
    x"CD",x"69",x"0D",x"F1",x"FC",x"20",x"0D",x"AF", -- 0x0B90
    x"32",x"1C",x"41",x"F1",x"D0",x"C3",x"D8",x"0C", -- 0x0B98
    x"21",x"1D",x"41",x"7E",x"35",x"B7",x"23",x"28", -- 0x0BA0
    x"FA",x"C9",x"E5",x"21",x"00",x"00",x"78",x"B1", -- 0x0BA8
    x"28",x"12",x"3E",x"10",x"29",x"DA",x"3D",x"27", -- 0x0BB0
    x"EB",x"29",x"EB",x"30",x"04",x"09",x"DA",x"3D", -- 0x0BB8
    x"27",x"3D",x"20",x"F0",x"EB",x"E1",x"C9",x"7C", -- 0x0BC0
    x"17",x"9F",x"47",x"CD",x"51",x"0C",x"79",x"98", -- 0x0BC8
    x"18",x"03",x"7C",x"17",x"9F",x"47",x"E5",x"7A", -- 0x0BD0
    x"17",x"9F",x"19",x"88",x"0F",x"AC",x"F2",x"99", -- 0x0BD8
    x"0A",x"C5",x"EB",x"CD",x"CF",x"0A",x"F1",x"E1", -- 0x0BE0
    x"CD",x"A4",x"09",x"EB",x"CD",x"6B",x"0C",x"C3", -- 0x0BE8
    x"8F",x"0F",x"7C",x"B5",x"CA",x"9A",x"0A",x"E5", -- 0x0BF0
    x"D5",x"CD",x"45",x"0C",x"C5",x"44",x"4D",x"21", -- 0x0BF8
    x"00",x"00",x"3E",x"10",x"29",x"38",x"1F",x"EB", -- 0x0C00
    x"29",x"EB",x"30",x"04",x"09",x"DA",x"26",x"0C", -- 0x0C08
    x"3D",x"20",x"F1",x"C1",x"D1",x"7C",x"B7",x"FA", -- 0x0C10
    x"1F",x"0C",x"D1",x"78",x"C3",x"4D",x"0C",x"EE", -- 0x0C18
    x"80",x"B5",x"28",x"13",x"EB",x"01",x"C1",x"E1", -- 0x0C20
    x"CD",x"CF",x"0A",x"E1",x"CD",x"A4",x"09",x"CD", -- 0x0C28
    x"CF",x"0A",x"C1",x"D1",x"C3",x"47",x"08",x"78", -- 0x0C30
    x"B7",x"C1",x"FA",x"9A",x"0A",x"D5",x"CD",x"CF", -- 0x0C38
    x"0A",x"D1",x"C3",x"82",x"09",x"7C",x"AA",x"47", -- 0x0C40
    x"CD",x"4C",x"0C",x"EB",x"7C",x"B7",x"F2",x"9A", -- 0x0C48
    x"0A",x"AF",x"4F",x"95",x"6F",x"79",x"9C",x"67", -- 0x0C50
    x"C3",x"9A",x"0A",x"2A",x"21",x"41",x"CD",x"51", -- 0x0C58
    x"0C",x"7C",x"EE",x"80",x"B5",x"C0",x"EB",x"CD", -- 0x0C60
    x"EF",x"0A",x"AF",x"06",x"98",x"C3",x"69",x"09", -- 0x0C68
    x"21",x"2D",x"41",x"7E",x"EE",x"80",x"77",x"21", -- 0x0C70
    x"2E",x"41",x"7E",x"B7",x"C8",x"47",x"2B",x"4E", -- 0x0C78
    x"11",x"24",x"41",x"1A",x"B7",x"CA",x"F4",x"09", -- 0x0C80
    x"90",x"30",x"16",x"2F",x"3C",x"F5",x"0E",x"08", -- 0x0C88
    x"23",x"E5",x"1A",x"46",x"77",x"78",x"12",x"1B", -- 0x0C90
    x"2B",x"0D",x"20",x"F6",x"E1",x"46",x"2B",x"4E", -- 0x0C98
    x"F1",x"FE",x"39",x"D0",x"F5",x"CD",x"DF",x"09", -- 0x0CA0
    x"23",x"36",x"00",x"47",x"F1",x"21",x"2D",x"41", -- 0x0CA8
    x"CD",x"69",x"0D",x"3A",x"26",x"41",x"32",x"1C", -- 0x0CB0
    x"41",x"78",x"B7",x"F2",x"CF",x"0C",x"CD",x"33", -- 0x0CB8
    x"0D",x"D2",x"0E",x"0D",x"EB",x"34",x"CA",x"B2", -- 0x0CC0
    x"07",x"CD",x"90",x"0D",x"C3",x"0E",x"0D",x"CD", -- 0x0CC8
    x"45",x"0D",x"21",x"25",x"41",x"DC",x"57",x"0D", -- 0x0CD0
    x"AF",x"47",x"3A",x"23",x"41",x"B7",x"20",x"1E", -- 0x0CD8
    x"21",x"1C",x"41",x"0E",x"08",x"56",x"77",x"7A", -- 0x0CE0
    x"23",x"0D",x"20",x"F9",x"78",x"D6",x"08",x"FE", -- 0x0CE8
    x"C0",x"20",x"E6",x"C3",x"78",x"07",x"05",x"21", -- 0x0CF0
    x"1C",x"41",x"CD",x"97",x"0D",x"B7",x"F2",x"F6", -- 0x0CF8
    x"0C",x"78",x"B7",x"28",x"09",x"21",x"24",x"41", -- 0x0D00
    x"86",x"77",x"D2",x"78",x"07",x"C8",x"3A",x"1C", -- 0x0D08
    x"41",x"B7",x"FC",x"20",x"0D",x"21",x"25",x"41", -- 0x0D10
    x"7E",x"E6",x"80",x"2B",x"2B",x"AE",x"77",x"C9", -- 0x0D18
    x"21",x"1D",x"41",x"06",x"07",x"34",x"C0",x"23", -- 0x0D20
    x"05",x"20",x"FA",x"34",x"CA",x"B2",x"07",x"2B", -- 0x0D28
    x"36",x"80",x"C9",x"21",x"27",x"41",x"11",x"1D", -- 0x0D30
    x"41",x"0E",x"07",x"AF",x"1A",x"8E",x"12",x"13", -- 0x0D38
    x"23",x"0D",x"20",x"F8",x"C9",x"21",x"27",x"41", -- 0x0D40
    x"11",x"1D",x"41",x"0E",x"07",x"AF",x"1A",x"9E", -- 0x0D48
    x"12",x"13",x"23",x"0D",x"20",x"F8",x"C9",x"7E", -- 0x0D50
    x"2F",x"77",x"21",x"1C",x"41",x"06",x"08",x"AF", -- 0x0D58
    x"4F",x"79",x"9E",x"77",x"23",x"05",x"20",x"F9", -- 0x0D60
    x"C9",x"71",x"E5",x"D6",x"08",x"38",x"0E",x"E1", -- 0x0D68
    x"E5",x"11",x"00",x"08",x"4E",x"73",x"59",x"2B", -- 0x0D70
    x"15",x"20",x"F9",x"18",x"EE",x"C6",x"09",x"57", -- 0x0D78
    x"AF",x"E1",x"15",x"C8",x"E5",x"1E",x"08",x"7E", -- 0x0D80
    x"1F",x"77",x"2B",x"1D",x"20",x"F9",x"18",x"F0", -- 0x0D88
    x"21",x"23",x"41",x"16",x"01",x"18",x"ED",x"0E", -- 0x0D90
    x"08",x"7E",x"17",x"77",x"23",x"0D",x"20",x"F9", -- 0x0D98
    x"C9",x"CD",x"55",x"09",x"C8",x"CD",x"0A",x"09", -- 0x0DA0
    x"CD",x"39",x"0E",x"71",x"13",x"06",x"07",x"1A", -- 0x0DA8
    x"13",x"B7",x"D5",x"28",x"17",x"0E",x"08",x"C5", -- 0x0DB0
    x"1F",x"47",x"DC",x"33",x"0D",x"CD",x"90",x"0D", -- 0x0DB8
    x"78",x"C1",x"0D",x"20",x"F2",x"D1",x"05",x"20", -- 0x0DC0
    x"E6",x"C3",x"D8",x"0C",x"21",x"23",x"41",x"CD", -- 0x0DC8
    x"70",x"0D",x"18",x"F1",x"00",x"00",x"00",x"00", -- 0x0DD0
    x"00",x"00",x"20",x"84",x"11",x"D4",x"0D",x"21", -- 0x0DD8
    x"27",x"41",x"CD",x"D3",x"09",x"3A",x"2E",x"41", -- 0x0DE0
    x"B7",x"CA",x"9A",x"19",x"CD",x"07",x"09",x"34", -- 0x0DE8
    x"34",x"CD",x"39",x"0E",x"21",x"51",x"41",x"71", -- 0x0DF0
    x"41",x"11",x"4A",x"41",x"21",x"27",x"41",x"CD", -- 0x0DF8
    x"4B",x"0D",x"1A",x"99",x"3F",x"38",x"0B",x"11", -- 0x0E00
    x"4A",x"41",x"21",x"27",x"41",x"CD",x"39",x"0D", -- 0x0E08
    x"AF",x"DA",x"12",x"04",x"3A",x"23",x"41",x"3C", -- 0x0E10
    x"3D",x"1F",x"FA",x"11",x"0D",x"17",x"21",x"1D", -- 0x0E18
    x"41",x"0E",x"07",x"CD",x"99",x"0D",x"21",x"4A", -- 0x0E20
    x"41",x"CD",x"97",x"0D",x"78",x"B7",x"20",x"C9", -- 0x0E28
    x"21",x"24",x"41",x"35",x"20",x"C3",x"C3",x"B2", -- 0x0E30
    x"07",x"79",x"32",x"2D",x"41",x"2B",x"11",x"50", -- 0x0E38
    x"41",x"01",x"00",x"07",x"7E",x"12",x"71",x"1B", -- 0x0E40
    x"2B",x"05",x"20",x"F8",x"C9",x"CD",x"FC",x"09", -- 0x0E48
    x"EB",x"2B",x"7E",x"B7",x"C8",x"C6",x"02",x"DA", -- 0x0E50
    x"B2",x"07",x"77",x"E5",x"CD",x"77",x"0C",x"E1", -- 0x0E58
    x"34",x"C0",x"C3",x"B2",x"07",x"CD",x"78",x"07", -- 0x0E60
    x"CD",x"EC",x"0A",x"F6",x"AF",x"EB",x"01",x"FF", -- 0x0E68
    x"00",x"60",x"68",x"CC",x"9A",x"0A",x"EB",x"7E", -- 0x0E70
    x"FE",x"2D",x"F5",x"CA",x"83",x"0E",x"FE",x"2B", -- 0x0E78
    x"28",x"01",x"2B",x"D7",x"DA",x"29",x"0F",x"FE", -- 0x0E80
    x"2E",x"CA",x"E4",x"0E",x"FE",x"45",x"28",x"14", -- 0x0E88
    x"FE",x"25",x"CA",x"EE",x"0E",x"FE",x"23",x"CA", -- 0x0E90
    x"F5",x"0E",x"FE",x"21",x"CA",x"F6",x"0E",x"FE", -- 0x0E98
    x"44",x"20",x"24",x"B7",x"CD",x"FB",x"0E",x"E5", -- 0x0EA0
    x"21",x"BD",x"0E",x"E3",x"D7",x"15",x"FE",x"CE", -- 0x0EA8
    x"C8",x"FE",x"2D",x"C8",x"14",x"FE",x"CD",x"C8", -- 0x0EB0
    x"FE",x"2B",x"C8",x"2B",x"F1",x"D7",x"DA",x"94", -- 0x0EB8
    x"0F",x"14",x"20",x"03",x"AF",x"93",x"5F",x"E5", -- 0x0EC0
    x"7B",x"90",x"F4",x"0A",x"0F",x"FC",x"18",x"0F", -- 0x0EC8
    x"20",x"F8",x"E1",x"F1",x"E5",x"CC",x"7B",x"09", -- 0x0ED0
    x"E1",x"E7",x"E8",x"E5",x"21",x"90",x"08",x"E5", -- 0x0ED8
    x"CD",x"A3",x"0A",x"C9",x"E7",x"0C",x"20",x"DF", -- 0x0EE0
    x"DC",x"FB",x"0E",x"C3",x"83",x"0E",x"E7",x"F2", -- 0x0EE8
    x"97",x"19",x"23",x"18",x"D2",x"B7",x"CD",x"FB", -- 0x0EF0
    x"0E",x"18",x"F7",x"E5",x"D5",x"C5",x"F5",x"CC", -- 0x0EF8
    x"B1",x"0A",x"F1",x"C4",x"DB",x"0A",x"C1",x"D1", -- 0x0F00
    x"E1",x"C9",x"C8",x"F5",x"E7",x"F5",x"E4",x"3E", -- 0x0F08
    x"09",x"F1",x"EC",x"4D",x"0E",x"F1",x"3D",x"C9", -- 0x0F10
    x"D5",x"E5",x"F5",x"E7",x"F5",x"E4",x"97",x"08", -- 0x0F18
    x"F1",x"EC",x"DC",x"0D",x"F1",x"E1",x"D1",x"3C", -- 0x0F20
    x"C9",x"D5",x"78",x"89",x"47",x"C5",x"E5",x"7E", -- 0x0F28
    x"D6",x"30",x"F5",x"E7",x"F2",x"5D",x"0F",x"2A", -- 0x0F30
    x"21",x"41",x"11",x"CD",x"0C",x"DF",x"30",x"19", -- 0x0F38
    x"54",x"5D",x"29",x"29",x"19",x"29",x"F1",x"4F", -- 0x0F40
    x"09",x"7C",x"B7",x"FA",x"57",x"0F",x"22",x"21", -- 0x0F48
    x"41",x"E1",x"C1",x"D1",x"C3",x"83",x"0E",x"79", -- 0x0F50
    x"F5",x"CD",x"CC",x"0A",x"37",x"30",x"18",x"01", -- 0x0F58
    x"74",x"94",x"11",x"00",x"24",x"CD",x"0C",x"0A", -- 0x0F60
    x"F2",x"74",x"0F",x"CD",x"3E",x"09",x"F1",x"CD", -- 0x0F68
    x"89",x"0F",x"18",x"DD",x"CD",x"E3",x"0A",x"CD", -- 0x0F70
    x"4D",x"0E",x"CD",x"FC",x"09",x"F1",x"CD",x"64", -- 0x0F78
    x"09",x"CD",x"E3",x"0A",x"CD",x"77",x"0C",x"18", -- 0x0F80
    x"C8",x"CD",x"A4",x"09",x"CD",x"64",x"09",x"C1", -- 0x0F88
    x"D1",x"C3",x"16",x"07",x"7B",x"FE",x"0A",x"30", -- 0x0F90
    x"09",x"07",x"07",x"83",x"07",x"86",x"D6",x"30", -- 0x0F98
    x"5F",x"FA",x"1E",x"32",x"C3",x"BD",x"0E",x"E5", -- 0x0FA0
    x"21",x"24",x"19",x"CD",x"A7",x"28",x"E1",x"CD", -- 0x0FA8
    x"9A",x"0A",x"AF",x"CD",x"34",x"10",x"B6",x"CD", -- 0x0FB0
    x"D9",x"0F",x"C3",x"A6",x"28",x"AF",x"CD",x"34", -- 0x0FB8
    x"10",x"E6",x"08",x"28",x"02",x"36",x"2B",x"EB", -- 0x0FC0
    x"CD",x"94",x"09",x"EB",x"F2",x"D9",x"0F",x"36", -- 0x0FC8
    x"2D",x"C5",x"E5",x"CD",x"7B",x"09",x"E1",x"C1", -- 0x0FD0
    x"B4",x"23",x"36",x"30",x"3A",x"D8",x"40",x"57", -- 0x0FD8
    x"17",x"3A",x"AF",x"40",x"DA",x"9A",x"10",x"CA", -- 0x0FE0
    x"92",x"10",x"FE",x"04",x"D2",x"3D",x"10",x"01", -- 0x0FE8
    x"00",x"00",x"CD",x"2F",x"13",x"21",x"30",x"41", -- 0x0FF0
    x"46",x"0E",x"20",x"3A",x"D8",x"40",x"5F",x"E6", -- 0x0FF8
    x"20",x"28",x"07",x"78",x"B9",x"0E",x"2A",x"20", -- 0x1000
    x"01",x"41",x"71",x"D7",x"28",x"14",x"FE",x"45", -- 0x1008
    x"28",x"10",x"FE",x"44",x"28",x"0C",x"FE",x"30", -- 0x1010
    x"28",x"F0",x"FE",x"2C",x"28",x"EC",x"FE",x"2E", -- 0x1018
    x"20",x"03",x"2B",x"36",x"30",x"7B",x"E6",x"10", -- 0x1020
    x"28",x"03",x"2B",x"36",x"24",x"7B",x"E6",x"04", -- 0x1028
    x"C0",x"2B",x"70",x"C9",x"32",x"D8",x"40",x"21", -- 0x1030
    x"30",x"41",x"36",x"20",x"C9",x"FE",x"05",x"E5", -- 0x1038
    x"DE",x"00",x"17",x"57",x"14",x"CD",x"01",x"12", -- 0x1040
    x"01",x"00",x"03",x"82",x"FA",x"57",x"10",x"14", -- 0x1048
    x"BA",x"30",x"04",x"3C",x"47",x"3E",x"02",x"D6", -- 0x1050
    x"02",x"E1",x"F5",x"CD",x"91",x"12",x"36",x"30", -- 0x1058
    x"CC",x"C9",x"09",x"CD",x"A4",x"12",x"2B",x"7E", -- 0x1060
    x"FE",x"30",x"28",x"FA",x"FE",x"2E",x"C4",x"C9", -- 0x1068
    x"09",x"F1",x"28",x"1F",x"F5",x"E7",x"3E",x"22", -- 0x1070
    x"8F",x"77",x"23",x"F1",x"36",x"2B",x"F2",x"85", -- 0x1078
    x"10",x"36",x"2D",x"2F",x"3C",x"06",x"2F",x"04", -- 0x1080
    x"D6",x"0A",x"30",x"FB",x"C6",x"3A",x"23",x"70", -- 0x1088
    x"23",x"77",x"23",x"36",x"00",x"EB",x"21",x"30", -- 0x1090
    x"41",x"C9",x"23",x"C5",x"FE",x"04",x"7A",x"D2", -- 0x1098
    x"09",x"11",x"1F",x"DA",x"A3",x"11",x"01",x"03", -- 0x10A0
    x"06",x"CD",x"89",x"12",x"D1",x"7A",x"D6",x"05", -- 0x10A8
    x"F4",x"69",x"12",x"CD",x"2F",x"13",x"7B",x"B7", -- 0x10B0
    x"CC",x"2F",x"09",x"3D",x"F4",x"69",x"12",x"E5", -- 0x10B8
    x"CD",x"F5",x"0F",x"E1",x"28",x"02",x"70",x"23", -- 0x10C0
    x"36",x"00",x"21",x"2F",x"41",x"23",x"3A",x"F3", -- 0x10C8
    x"40",x"95",x"92",x"C8",x"7E",x"FE",x"20",x"28", -- 0x10D0
    x"F4",x"FE",x"2A",x"28",x"F0",x"2B",x"E5",x"F5", -- 0x10D8
    x"01",x"DF",x"10",x"C5",x"D7",x"FE",x"2D",x"C8", -- 0x10E0
    x"FE",x"2B",x"C8",x"FE",x"24",x"C8",x"C1",x"FE", -- 0x10E8
    x"30",x"20",x"0F",x"23",x"D7",x"30",x"0B",x"2B", -- 0x10F0
    x"01",x"2B",x"77",x"F1",x"28",x"FB",x"C1",x"C3", -- 0x10F8
    x"CE",x"10",x"F1",x"28",x"FD",x"E1",x"36",x"25", -- 0x1100
    x"C9",x"E5",x"1F",x"DA",x"AA",x"11",x"28",x"14", -- 0x1108
    x"11",x"84",x"13",x"CD",x"49",x"0A",x"16",x"10", -- 0x1110
    x"FA",x"32",x"11",x"E1",x"C1",x"CD",x"BD",x"0F", -- 0x1118
    x"2B",x"36",x"25",x"C9",x"01",x"0E",x"B6",x"11", -- 0x1120
    x"CA",x"1B",x"CD",x"0C",x"0A",x"F2",x"1B",x"11", -- 0x1128
    x"16",x"06",x"CD",x"55",x"09",x"C4",x"01",x"12", -- 0x1130
    x"E1",x"C1",x"FA",x"57",x"11",x"C5",x"5F",x"78", -- 0x1138
    x"92",x"93",x"F4",x"69",x"12",x"CD",x"7D",x"12", -- 0x1140
    x"CD",x"A4",x"12",x"B3",x"C4",x"77",x"12",x"B3", -- 0x1148
    x"C4",x"91",x"12",x"D1",x"C3",x"B6",x"10",x"5F", -- 0x1150
    x"79",x"B7",x"C4",x"16",x"0F",x"83",x"FA",x"62", -- 0x1158
    x"11",x"AF",x"C5",x"F5",x"FC",x"18",x"0F",x"FA", -- 0x1160
    x"64",x"11",x"C1",x"7B",x"90",x"C1",x"5F",x"82", -- 0x1168
    x"78",x"FA",x"7F",x"11",x"92",x"93",x"F4",x"69", -- 0x1170
    x"12",x"C5",x"CD",x"7D",x"12",x"18",x"11",x"CD", -- 0x1178
    x"69",x"12",x"79",x"CD",x"94",x"12",x"4F",x"AF", -- 0x1180
    x"92",x"93",x"CD",x"69",x"12",x"C5",x"47",x"4F", -- 0x1188
    x"CD",x"A4",x"12",x"C1",x"B1",x"20",x"03",x"2A", -- 0x1190
    x"F3",x"40",x"83",x"3D",x"F4",x"69",x"12",x"50", -- 0x1198
    x"C3",x"BF",x"10",x"E5",x"D5",x"CD",x"CC",x"0A", -- 0x11A0
    x"D1",x"AF",x"CA",x"B0",x"11",x"1E",x"10",x"01", -- 0x11A8
    x"1E",x"06",x"CD",x"55",x"09",x"37",x"C4",x"01", -- 0x11B0
    x"12",x"E1",x"C1",x"F5",x"79",x"B7",x"F5",x"C4", -- 0x11B8
    x"16",x"0F",x"80",x"4F",x"7A",x"E6",x"04",x"FE", -- 0x11C0
    x"01",x"9F",x"57",x"81",x"4F",x"93",x"F5",x"C5", -- 0x11C8
    x"FC",x"18",x"0F",x"FA",x"D0",x"11",x"C1",x"F1", -- 0x11D0
    x"C5",x"F5",x"FA",x"DE",x"11",x"AF",x"2F",x"3C", -- 0x11D8
    x"80",x"3C",x"82",x"47",x"0E",x"00",x"CD",x"A4", -- 0x11E0
    x"12",x"F1",x"F4",x"71",x"12",x"C1",x"F1",x"CC", -- 0x11E8
    x"2F",x"09",x"F1",x"38",x"03",x"83",x"90",x"92", -- 0x11F0
    x"C5",x"CD",x"74",x"10",x"EB",x"D1",x"C3",x"BF", -- 0x11F8
    x"10",x"D5",x"AF",x"F5",x"E7",x"E2",x"22",x"12", -- 0x1200
    x"3A",x"24",x"41",x"FE",x"91",x"D2",x"22",x"12", -- 0x1208
    x"11",x"64",x"13",x"21",x"27",x"41",x"CD",x"D3", -- 0x1210
    x"09",x"CD",x"A1",x"0D",x"F1",x"D6",x"0A",x"F5", -- 0x1218
    x"18",x"E6",x"CD",x"4F",x"12",x"E7",x"30",x"0B", -- 0x1220
    x"01",x"43",x"91",x"11",x"F9",x"4F",x"CD",x"0C", -- 0x1228
    x"0A",x"18",x"06",x"11",x"6C",x"13",x"CD",x"49", -- 0x1230
    x"0A",x"F2",x"4B",x"12",x"F1",x"CD",x"0B",x"0F", -- 0x1238
    x"F5",x"18",x"E2",x"F1",x"CD",x"18",x"0F",x"F5", -- 0x1240
    x"CD",x"4F",x"12",x"F1",x"B7",x"D1",x"C9",x"E7", -- 0x1248
    x"EA",x"5E",x"12",x"01",x"74",x"94",x"11",x"F8", -- 0x1250
    x"23",x"CD",x"0C",x"0A",x"18",x"06",x"11",x"74", -- 0x1258
    x"13",x"CD",x"49",x"0A",x"E1",x"F2",x"43",x"12", -- 0x1260
    x"E9",x"B7",x"C8",x"3D",x"36",x"30",x"23",x"18", -- 0x1268
    x"F9",x"20",x"04",x"C8",x"CD",x"91",x"12",x"36", -- 0x1270
    x"30",x"23",x"3D",x"18",x"F6",x"7B",x"82",x"3C", -- 0x1278
    x"47",x"3C",x"D6",x"03",x"30",x"FC",x"C6",x"05", -- 0x1280
    x"4F",x"3A",x"D8",x"40",x"E6",x"40",x"C0",x"4F", -- 0x1288
    x"C9",x"05",x"20",x"08",x"36",x"2E",x"22",x"F3", -- 0x1290
    x"40",x"23",x"48",x"C9",x"0D",x"C0",x"36",x"2C", -- 0x1298
    x"23",x"0E",x"03",x"C9",x"D5",x"E7",x"E2",x"EA", -- 0x12A0
    x"12",x"C5",x"E5",x"CD",x"FC",x"09",x"21",x"7C", -- 0x12A8
    x"13",x"CD",x"F7",x"09",x"CD",x"77",x"0C",x"AF", -- 0x12B0
    x"CD",x"7B",x"0B",x"E1",x"C1",x"11",x"8C",x"13", -- 0x12B8
    x"3E",x"0A",x"CD",x"91",x"12",x"C5",x"F5",x"E5", -- 0x12C0
    x"D5",x"06",x"2F",x"04",x"E1",x"E5",x"CD",x"48", -- 0x12C8
    x"0D",x"30",x"F8",x"E1",x"CD",x"36",x"0D",x"EB", -- 0x12D0
    x"E1",x"70",x"23",x"F1",x"C1",x"3D",x"20",x"E2", -- 0x12D8
    x"C5",x"E5",x"21",x"1D",x"41",x"CD",x"B1",x"09", -- 0x12E0
    x"18",x"0C",x"C5",x"E5",x"CD",x"08",x"07",x"3C", -- 0x12E8
    x"CD",x"FB",x"0A",x"CD",x"B4",x"09",x"E1",x"C1", -- 0x12F0
    x"AF",x"11",x"D2",x"13",x"3F",x"CD",x"91",x"12", -- 0x12F8
    x"C5",x"F5",x"E5",x"D5",x"CD",x"BF",x"09",x"E1", -- 0x1300
    x"06",x"2F",x"04",x"7B",x"96",x"5F",x"23",x"7A", -- 0x1308
    x"9E",x"57",x"23",x"79",x"9E",x"4F",x"2B",x"2B", -- 0x1310
    x"30",x"F0",x"CD",x"B7",x"07",x"23",x"CD",x"B4", -- 0x1318
    x"09",x"EB",x"E1",x"70",x"23",x"F1",x"C1",x"38", -- 0x1320
    x"D3",x"13",x"13",x"3E",x"04",x"18",x"06",x"D5", -- 0x1328
    x"11",x"D8",x"13",x"3E",x"05",x"CD",x"91",x"12", -- 0x1330
    x"C5",x"F5",x"E5",x"EB",x"4E",x"23",x"46",x"C5", -- 0x1338
    x"23",x"E3",x"EB",x"2A",x"21",x"41",x"06",x"2F", -- 0x1340
    x"04",x"7D",x"93",x"6F",x"7C",x"9A",x"67",x"30", -- 0x1348
    x"F7",x"19",x"22",x"21",x"41",x"D1",x"E1",x"70", -- 0x1350
    x"23",x"F1",x"C1",x"3D",x"20",x"D7",x"CD",x"91", -- 0x1358
    x"12",x"77",x"D1",x"C9",x"00",x"00",x"00",x"00", -- 0x1360
    x"F9",x"02",x"15",x"A2",x"FD",x"FF",x"9F",x"31", -- 0x1368
    x"A9",x"5F",x"63",x"B2",x"FE",x"FF",x"03",x"BF", -- 0x1370
    x"C9",x"1B",x"0E",x"B6",x"00",x"00",x"00",x"00", -- 0x1378
    x"00",x"00",x"00",x"80",x"00",x"00",x"04",x"BF", -- 0x1380
    x"C9",x"1B",x"0E",x"B6",x"00",x"80",x"C6",x"A4", -- 0x1388
    x"7E",x"8D",x"03",x"00",x"40",x"7A",x"10",x"F3", -- 0x1390
    x"5A",x"00",x"00",x"A0",x"72",x"4E",x"18",x"09", -- 0x1398
    x"00",x"00",x"10",x"A5",x"D4",x"E8",x"00",x"00", -- 0x13A0
    x"00",x"E8",x"76",x"48",x"17",x"00",x"00",x"00", -- 0x13A8
    x"E4",x"0B",x"54",x"02",x"00",x"00",x"00",x"CA", -- 0x13B0
    x"9A",x"3B",x"00",x"00",x"00",x"00",x"E1",x"F5", -- 0x13B8
    x"05",x"00",x"00",x"00",x"80",x"96",x"98",x"00", -- 0x13C0
    x"00",x"00",x"00",x"40",x"42",x"0F",x"00",x"00", -- 0x13C8
    x"00",x"00",x"A0",x"86",x"01",x"10",x"27",x"00", -- 0x13D0
    x"10",x"27",x"E8",x"03",x"64",x"00",x"0A",x"00", -- 0x13D8
    x"01",x"00",x"21",x"82",x"09",x"E3",x"E9",x"CD", -- 0x13E0
    x"A4",x"09",x"21",x"80",x"13",x"CD",x"B1",x"09", -- 0x13E8
    x"18",x"03",x"CD",x"B1",x"0A",x"C1",x"D1",x"CD", -- 0x13F0
    x"55",x"09",x"78",x"28",x"3C",x"F2",x"04",x"14", -- 0x13F8
    x"B7",x"CA",x"9A",x"19",x"B7",x"CA",x"79",x"07", -- 0x1400
    x"D5",x"C5",x"79",x"F6",x"7F",x"CD",x"BF",x"09", -- 0x1408
    x"F2",x"21",x"14",x"D5",x"C5",x"CD",x"40",x"0B", -- 0x1410
    x"C1",x"D1",x"F5",x"CD",x"0C",x"0A",x"E1",x"7C", -- 0x1418
    x"1F",x"E1",x"22",x"23",x"41",x"E1",x"22",x"21", -- 0x1420
    x"41",x"DC",x"E2",x"13",x"CC",x"82",x"09",x"D5", -- 0x1428
    x"C5",x"CD",x"09",x"08",x"C1",x"D1",x"CD",x"47", -- 0x1430
    x"08",x"CD",x"A4",x"09",x"01",x"38",x"81",x"11", -- 0x1438
    x"3B",x"AA",x"CD",x"47",x"08",x"3A",x"24",x"41", -- 0x1440
    x"FE",x"88",x"D2",x"31",x"09",x"CD",x"40",x"0B", -- 0x1448
    x"C6",x"80",x"C6",x"02",x"DA",x"31",x"09",x"F5", -- 0x1450
    x"21",x"F8",x"07",x"CD",x"0B",x"07",x"CD",x"41", -- 0x1458
    x"08",x"F1",x"C1",x"D1",x"F5",x"CD",x"13",x"07", -- 0x1460
    x"CD",x"82",x"09",x"21",x"79",x"14",x"CD",x"A9", -- 0x1468
    x"14",x"11",x"00",x"00",x"C1",x"4A",x"C3",x"47", -- 0x1470
    x"08",x"08",x"40",x"2E",x"94",x"74",x"70",x"4F", -- 0x1478
    x"2E",x"77",x"6E",x"02",x"88",x"7A",x"E6",x"A0", -- 0x1480
    x"2A",x"7C",x"50",x"AA",x"AA",x"7E",x"FF",x"FF", -- 0x1488
    x"7F",x"7F",x"00",x"00",x"80",x"81",x"00",x"00", -- 0x1490
    x"00",x"81",x"CD",x"A4",x"09",x"11",x"32",x"0C", -- 0x1498
    x"D5",x"E5",x"CD",x"BF",x"09",x"CD",x"47",x"08", -- 0x14A0
    x"E1",x"CD",x"A4",x"09",x"7E",x"23",x"CD",x"B1", -- 0x14A8
    x"09",x"06",x"F1",x"C1",x"D1",x"3D",x"C8",x"D5", -- 0x14B0
    x"C5",x"F5",x"E5",x"CD",x"47",x"08",x"E1",x"CD", -- 0x14B8
    x"C2",x"09",x"E5",x"CD",x"16",x"07",x"E1",x"18", -- 0x14C0
    x"E9",x"CD",x"7F",x"0A",x"7C",x"B7",x"FA",x"4A", -- 0x14C8
    x"1E",x"B5",x"CA",x"F0",x"14",x"E5",x"CD",x"F0", -- 0x14D0
    x"14",x"CD",x"BF",x"09",x"EB",x"E3",x"C5",x"CD", -- 0x14D8
    x"CF",x"0A",x"C1",x"D1",x"CD",x"47",x"08",x"21", -- 0x14E0
    x"F8",x"07",x"CD",x"0B",x"07",x"C3",x"40",x"0B", -- 0x14E8
    x"21",x"90",x"40",x"E5",x"11",x"00",x"00",x"4B", -- 0x14F0
    x"26",x"03",x"2E",x"08",x"EB",x"29",x"EB",x"79", -- 0x14F8
    x"17",x"4F",x"E3",x"7E",x"07",x"77",x"E3",x"D2", -- 0x1500
    x"16",x"15",x"E5",x"2A",x"AA",x"40",x"19",x"EB", -- 0x1508
    x"3A",x"AC",x"40",x"89",x"4F",x"E1",x"2D",x"C2", -- 0x1510
    x"FC",x"14",x"E3",x"23",x"E3",x"25",x"C2",x"FA", -- 0x1518
    x"14",x"E1",x"21",x"65",x"B0",x"19",x"22",x"AA", -- 0x1520
    x"40",x"CD",x"EF",x"0A",x"3E",x"05",x"89",x"32", -- 0x1528
    x"AC",x"40",x"EB",x"06",x"80",x"21",x"25",x"41", -- 0x1530
    x"70",x"2B",x"70",x"4F",x"06",x"00",x"C3",x"65", -- 0x1538
    x"07",x"21",x"8B",x"15",x"CD",x"0B",x"07",x"CD", -- 0x1540
    x"A4",x"09",x"01",x"49",x"83",x"11",x"DB",x"0F", -- 0x1548
    x"CD",x"B4",x"09",x"C1",x"D1",x"CD",x"A2",x"08", -- 0x1550
    x"CD",x"A4",x"09",x"CD",x"40",x"0B",x"C1",x"D1", -- 0x1558
    x"CD",x"13",x"07",x"21",x"8F",x"15",x"CD",x"10", -- 0x1560
    x"07",x"CD",x"55",x"09",x"37",x"F2",x"77",x"15", -- 0x1568
    x"CD",x"08",x"07",x"CD",x"55",x"09",x"B7",x"F5", -- 0x1570
    x"F4",x"82",x"09",x"21",x"8F",x"15",x"CD",x"0B", -- 0x1578
    x"07",x"F1",x"D4",x"82",x"09",x"21",x"93",x"15", -- 0x1580
    x"C3",x"9A",x"14",x"DB",x"0F",x"49",x"81",x"00", -- 0x1588
    x"00",x"00",x"7F",x"05",x"BA",x"D7",x"1E",x"86", -- 0x1590
    x"64",x"26",x"99",x"87",x"58",x"34",x"23",x"87", -- 0x1598
    x"E0",x"5D",x"A5",x"86",x"DA",x"0F",x"49",x"83", -- 0x15A0
    x"CD",x"A4",x"09",x"CD",x"47",x"15",x"C1",x"E1", -- 0x15A8
    x"CD",x"A4",x"09",x"EB",x"CD",x"B4",x"09",x"CD", -- 0x15B0
    x"41",x"15",x"C3",x"A0",x"08",x"CD",x"55",x"09", -- 0x15B8
    x"FC",x"E2",x"13",x"FC",x"82",x"09",x"3A",x"24", -- 0x15C0
    x"41",x"FE",x"81",x"38",x"0C",x"01",x"00",x"81", -- 0x15C8
    x"51",x"59",x"CD",x"A2",x"08",x"21",x"10",x"07", -- 0x15D0
    x"E5",x"21",x"E3",x"15",x"CD",x"9A",x"14",x"21", -- 0x15D8
    x"8B",x"15",x"C9",x"09",x"4A",x"D7",x"3B",x"78", -- 0x15E0
    x"02",x"6E",x"84",x"7B",x"FE",x"C1",x"2F",x"7C", -- 0x15E8
    x"74",x"31",x"9A",x"7D",x"84",x"3D",x"5A",x"7D", -- 0x15F0
    x"C8",x"7F",x"91",x"7E",x"E4",x"BB",x"4C",x"7E", -- 0x15F8
    x"6C",x"AA",x"AA",x"7F",x"00",x"00",x"00",x"81", -- 0x1600
    x"8A",x"09",x"37",x"0B",x"77",x"09",x"D4",x"27", -- 0x1608
    x"EF",x"2A",x"F5",x"27",x"E7",x"13",x"C9",x"14", -- 0x1610
    x"09",x"08",x"39",x"14",x"41",x"15",x"47",x"15", -- 0x1618
    x"A8",x"15",x"BD",x"15",x"AA",x"2C",x"52",x"41", -- 0x1620
    x"58",x"41",x"5E",x"41",x"61",x"41",x"64",x"41", -- 0x1628
    x"67",x"41",x"6A",x"41",x"6D",x"41",x"70",x"41", -- 0x1630
    x"7F",x"0A",x"B1",x"0A",x"DB",x"0A",x"26",x"0B", -- 0x1638
    x"03",x"2A",x"36",x"28",x"C5",x"2A",x"0F",x"2A", -- 0x1640
    x"1F",x"2A",x"61",x"2A",x"91",x"2A",x"9A",x"2A", -- 0x1648
    x"C5",x"4E",x"44",x"C6",x"4F",x"52",x"D2",x"45", -- 0x1650
    x"53",x"45",x"54",x"D3",x"45",x"54",x"C3",x"4C", -- 0x1658
    x"53",x"C3",x"4D",x"44",x"D2",x"41",x"4E",x"44", -- 0x1660
    x"4F",x"4D",x"CE",x"45",x"58",x"54",x"C4",x"41", -- 0x1668
    x"54",x"41",x"C9",x"4E",x"50",x"55",x"54",x"C4", -- 0x1670
    x"49",x"4D",x"D2",x"45",x"41",x"44",x"CC",x"45", -- 0x1678
    x"54",x"C7",x"4F",x"54",x"4F",x"D2",x"55",x"4E", -- 0x1680
    x"C9",x"46",x"D2",x"45",x"53",x"54",x"4F",x"52", -- 0x1688
    x"45",x"C7",x"4F",x"53",x"55",x"42",x"D2",x"45", -- 0x1690
    x"54",x"55",x"52",x"4E",x"D2",x"45",x"4D",x"D3", -- 0x1698
    x"54",x"4F",x"50",x"C5",x"4C",x"53",x"45",x"D4", -- 0x16A0
    x"52",x"4F",x"4E",x"D4",x"52",x"4F",x"46",x"46", -- 0x16A8
    x"C4",x"45",x"46",x"53",x"54",x"52",x"C4",x"45", -- 0x16B0
    x"46",x"49",x"4E",x"54",x"C4",x"45",x"46",x"53", -- 0x16B8
    x"4E",x"47",x"C4",x"45",x"46",x"44",x"42",x"4C", -- 0x16C0
    x"CC",x"49",x"4E",x"45",x"C5",x"44",x"49",x"54", -- 0x16C8
    x"C5",x"52",x"52",x"4F",x"52",x"D2",x"45",x"53", -- 0x16D0
    x"55",x"4D",x"45",x"CF",x"55",x"54",x"CF",x"4E", -- 0x16D8
    x"CF",x"50",x"45",x"4E",x"C6",x"49",x"45",x"4C", -- 0x16E0
    x"44",x"C7",x"45",x"54",x"D0",x"55",x"54",x"C3", -- 0x16E8
    x"4C",x"4F",x"53",x"45",x"CC",x"4F",x"41",x"44", -- 0x16F0
    x"CD",x"45",x"52",x"47",x"45",x"CE",x"41",x"4D", -- 0x16F8
    x"45",x"CB",x"49",x"4C",x"4C",x"CC",x"53",x"45", -- 0x1700
    x"54",x"D2",x"53",x"45",x"54",x"D3",x"41",x"56", -- 0x1708
    x"45",x"D3",x"59",x"53",x"54",x"45",x"4D",x"CC", -- 0x1710
    x"50",x"52",x"49",x"4E",x"54",x"C4",x"45",x"46", -- 0x1718
    x"D0",x"4F",x"4B",x"45",x"D0",x"52",x"49",x"4E", -- 0x1720
    x"54",x"C3",x"4F",x"4E",x"54",x"CC",x"49",x"53", -- 0x1728
    x"54",x"CC",x"4C",x"49",x"53",x"54",x"C4",x"45", -- 0x1730
    x"4C",x"45",x"54",x"45",x"C1",x"55",x"54",x"4F", -- 0x1738
    x"C3",x"4C",x"45",x"41",x"52",x"C3",x"4C",x"4F", -- 0x1740
    x"41",x"44",x"C3",x"53",x"41",x"56",x"45",x"CE", -- 0x1748
    x"45",x"57",x"D4",x"41",x"42",x"28",x"D4",x"4F", -- 0x1750
    x"C6",x"4E",x"D5",x"53",x"49",x"4E",x"47",x"D6", -- 0x1758
    x"41",x"52",x"50",x"54",x"52",x"D5",x"53",x"52", -- 0x1760
    x"C5",x"52",x"4C",x"C5",x"52",x"52",x"D3",x"54", -- 0x1768
    x"52",x"49",x"4E",x"47",x"24",x"C9",x"4E",x"53", -- 0x1770
    x"54",x"52",x"C3",x"48",x"45",x"43",x"4B",x"D4", -- 0x1778
    x"49",x"4D",x"45",x"24",x"CD",x"45",x"4D",x"C9", -- 0x1780
    x"4E",x"4B",x"45",x"59",x"24",x"D4",x"48",x"45", -- 0x1788
    x"4E",x"CE",x"4F",x"54",x"D3",x"54",x"45",x"50", -- 0x1790
    x"AB",x"AD",x"AA",x"AF",x"DB",x"C1",x"4E",x"44", -- 0x1798
    x"CF",x"52",x"BE",x"BD",x"BC",x"D3",x"47",x"4E", -- 0x17A0
    x"C9",x"4E",x"54",x"C1",x"42",x"53",x"C6",x"52", -- 0x17A8
    x"45",x"C9",x"4E",x"50",x"D0",x"4F",x"53",x"D3", -- 0x17B0
    x"51",x"52",x"D2",x"4E",x"44",x"CC",x"4F",x"47", -- 0x17B8
    x"C5",x"58",x"50",x"C3",x"4F",x"53",x"D3",x"49", -- 0x17C0
    x"4E",x"D4",x"41",x"4E",x"C1",x"54",x"4E",x"D0", -- 0x17C8
    x"45",x"45",x"4B",x"C3",x"56",x"49",x"C3",x"56", -- 0x17D0
    x"53",x"C3",x"56",x"44",x"C5",x"4F",x"46",x"CC", -- 0x17D8
    x"4F",x"43",x"CC",x"4F",x"46",x"CD",x"4B",x"49", -- 0x17E0
    x"24",x"CD",x"4B",x"53",x"24",x"CD",x"4B",x"44", -- 0x17E8
    x"24",x"C3",x"49",x"4E",x"54",x"C3",x"53",x"4E", -- 0x17F0
    x"47",x"C3",x"44",x"42",x"4C",x"C6",x"49",x"58", -- 0x17F8
    x"CC",x"45",x"4E",x"D3",x"54",x"52",x"24",x"D6", -- 0x1800
    x"41",x"4C",x"C1",x"53",x"43",x"C3",x"48",x"52", -- 0x1808
    x"24",x"CC",x"45",x"46",x"54",x"24",x"D2",x"49", -- 0x1810
    x"47",x"48",x"54",x"24",x"CD",x"49",x"44",x"24", -- 0x1818
    x"A7",x"80",x"AE",x"1D",x"A1",x"1C",x"38",x"01", -- 0x1820
    x"35",x"01",x"C9",x"01",x"73",x"41",x"D3",x"01", -- 0x1828
    x"B6",x"22",x"05",x"1F",x"9A",x"21",x"08",x"26", -- 0x1830
    x"EF",x"21",x"21",x"1F",x"C2",x"1E",x"A3",x"1E", -- 0x1838
    x"39",x"20",x"91",x"1D",x"B1",x"1E",x"DE",x"1E", -- 0x1840
    x"07",x"1F",x"A9",x"1D",x"07",x"1F",x"F7",x"1D", -- 0x1848
    x"F8",x"1D",x"00",x"1E",x"03",x"1E",x"06",x"1E", -- 0x1850
    x"09",x"1E",x"A3",x"41",x"60",x"2E",x"F4",x"1F", -- 0x1858
    x"AF",x"1F",x"FB",x"2A",x"6C",x"1F",x"79",x"41", -- 0x1860
    x"7C",x"41",x"7F",x"41",x"82",x"41",x"85",x"41", -- 0x1868
    x"88",x"41",x"8B",x"41",x"8E",x"41",x"91",x"41", -- 0x1870
    x"97",x"41",x"9A",x"41",x"A0",x"41",x"B2",x"02", -- 0x1878
    x"67",x"20",x"5B",x"41",x"B1",x"2C",x"6F",x"20", -- 0x1880
    x"E4",x"1D",x"2E",x"2B",x"29",x"2B",x"C6",x"2B", -- 0x1888
    x"08",x"20",x"7A",x"1E",x"1F",x"2C",x"F5",x"2B", -- 0x1890
    x"49",x"1B",x"79",x"79",x"7C",x"7C",x"7F",x"50", -- 0x1898
    x"46",x"DB",x"0A",x"00",x"00",x"7F",x"0A",x"F4", -- 0x18A0
    x"0A",x"B1",x"0A",x"77",x"0C",x"70",x"0C",x"A1", -- 0x18A8
    x"0D",x"E5",x"0D",x"78",x"0A",x"16",x"07",x"13", -- 0x18B0
    x"07",x"47",x"08",x"A2",x"08",x"0C",x"0A",x"D2", -- 0x18B8
    x"0B",x"C7",x"0B",x"F2",x"0B",x"90",x"24",x"39", -- 0x18C0
    x"0A",x"4E",x"46",x"53",x"4E",x"52",x"47",x"4F", -- 0x18C8
    x"44",x"46",x"43",x"4F",x"56",x"4F",x"4D",x"55", -- 0x18D0
    x"4C",x"42",x"53",x"44",x"44",x"2F",x"30",x"49", -- 0x18D8
    x"44",x"54",x"4D",x"4F",x"53",x"4C",x"53",x"53", -- 0x18E0
    x"54",x"43",x"4E",x"4E",x"52",x"52",x"57",x"55", -- 0x18E8
    x"45",x"4D",x"4F",x"46",x"44",x"53",x"4E",x"D6", -- 0x18F0
    x"00",x"6F",x"7C",x"DE",x"00",x"67",x"78",x"DE", -- 0x18F8
    x"00",x"47",x"3E",x"00",x"C9",x"4A",x"1E",x"40", -- 0x1900
    x"E6",x"4D",x"DB",x"00",x"C9",x"D3",x"00",x"C9", -- 0x1908
    x"00",x"00",x"00",x"00",x"28",x"1E",x"00",x"4C", -- 0x1910
    x"43",x"FE",x"FF",x"01",x"48",x"20",x"45",x"72", -- 0x1918
    x"72",x"6F",x"72",x"00",x"20",x"69",x"6E",x"20", -- 0x1920
    x"00",x"52",x"45",x"41",x"44",x"59",x"0D",x"00", -- 0x1928
    x"42",x"72",x"65",x"61",x"6B",x"00",x"21",x"04", -- 0x1930
    x"00",x"39",x"7E",x"23",x"FE",x"81",x"C0",x"4E", -- 0x1938
    x"23",x"46",x"23",x"E5",x"69",x"60",x"7A",x"B3", -- 0x1940
    x"EB",x"28",x"02",x"EB",x"DF",x"01",x"0E",x"00", -- 0x1948
    x"E1",x"C8",x"09",x"18",x"E5",x"CD",x"6C",x"19", -- 0x1950
    x"C5",x"E3",x"C1",x"DF",x"7E",x"02",x"C8",x"0B", -- 0x1958
    x"2B",x"18",x"F8",x"E5",x"2A",x"FD",x"40",x"06", -- 0x1960
    x"00",x"09",x"09",x"3E",x"E5",x"3E",x"C6",x"95", -- 0x1968
    x"6F",x"3E",x"FF",x"9C",x"38",x"04",x"67",x"39", -- 0x1970
    x"E1",x"D8",x"1E",x"0C",x"18",x"24",x"2A",x"A2", -- 0x1978
    x"40",x"7C",x"A5",x"3C",x"28",x"08",x"3A",x"F2", -- 0x1980
    x"40",x"B7",x"1E",x"22",x"20",x"14",x"C3",x"C1", -- 0x1988
    x"1D",x"2A",x"DA",x"40",x"22",x"A2",x"40",x"1E", -- 0x1990
    x"02",x"01",x"1E",x"14",x"01",x"1E",x"00",x"01", -- 0x1998
    x"1E",x"24",x"2A",x"A2",x"40",x"22",x"EA",x"40", -- 0x19A0
    x"22",x"EC",x"40",x"01",x"B4",x"19",x"2A",x"E8", -- 0x19A8
    x"40",x"C3",x"9A",x"1B",x"C1",x"7B",x"4B",x"32", -- 0x19B0
    x"9A",x"40",x"2A",x"E6",x"40",x"22",x"EE",x"40", -- 0x19B8
    x"EB",x"2A",x"EA",x"40",x"7C",x"A5",x"3C",x"28", -- 0x19C0
    x"07",x"22",x"F5",x"40",x"EB",x"22",x"F7",x"40", -- 0x19C8
    x"2A",x"F0",x"40",x"7C",x"B5",x"EB",x"21",x"F2", -- 0x19D0
    x"40",x"28",x"08",x"A6",x"20",x"05",x"35",x"EB", -- 0x19D8
    x"C3",x"36",x"1D",x"AF",x"77",x"59",x"CD",x"F9", -- 0x19E0
    x"20",x"21",x"C9",x"18",x"CD",x"A6",x"41",x"57", -- 0x19E8
    x"3E",x"3F",x"CD",x"2A",x"03",x"19",x"7E",x"CD", -- 0x19F0
    x"2A",x"03",x"D7",x"CD",x"2A",x"03",x"21",x"1D", -- 0x19F8
    x"19",x"E5",x"2A",x"EA",x"40",x"E3",x"CD",x"79", -- 0x1A00
    x"35",x"E1",x"11",x"FE",x"FF",x"DF",x"CA",x"74", -- 0x1A08
    x"06",x"7C",x"A5",x"3C",x"C4",x"A7",x"0F",x"3E", -- 0x1A10
    x"C1",x"CD",x"8B",x"03",x"CD",x"AC",x"41",x"00", -- 0x1A18
    x"00",x"00",x"CD",x"F9",x"20",x"21",x"29",x"19", -- 0x1A20
    x"CD",x"92",x"38",x"3A",x"9A",x"40",x"D6",x"02", -- 0x1A28
    x"CC",x"53",x"2E",x"21",x"FF",x"FF",x"22",x"A2", -- 0x1A30
    x"40",x"3A",x"E1",x"40",x"B7",x"28",x"37",x"2A", -- 0x1A38
    x"E2",x"40",x"E5",x"CD",x"AF",x"0F",x"D1",x"D5", -- 0x1A40
    x"CD",x"2C",x"1B",x"3E",x"2A",x"38",x"02",x"3E", -- 0x1A48
    x"20",x"CD",x"2A",x"03",x"CD",x"61",x"03",x"D1", -- 0x1A50
    x"30",x"06",x"AF",x"32",x"E1",x"40",x"18",x"B9", -- 0x1A58
    x"2A",x"E4",x"40",x"19",x"38",x"F4",x"D5",x"11", -- 0x1A60
    x"F9",x"FF",x"DF",x"D1",x"30",x"EC",x"22",x"E2", -- 0x1A68
    x"40",x"F6",x"FF",x"C3",x"EB",x"2F",x"3E",x"3E", -- 0x1A70
    x"CD",x"2A",x"03",x"CD",x"61",x"03",x"DA",x"33", -- 0x1A78
    x"1A",x"D7",x"3C",x"3D",x"CA",x"33",x"1A",x"F5", -- 0x1A80
    x"CD",x"5A",x"1E",x"2B",x"7E",x"FE",x"20",x"28", -- 0x1A88
    x"FA",x"23",x"7E",x"FE",x"20",x"CC",x"C9",x"09", -- 0x1A90
    x"D5",x"CD",x"C0",x"1B",x"D1",x"F1",x"22",x"E6", -- 0x1A98
    x"40",x"CD",x"B2",x"41",x"D2",x"5A",x"1D",x"D5", -- 0x1AA0
    x"C5",x"AF",x"32",x"DD",x"40",x"D7",x"B7",x"F5", -- 0x1AA8
    x"EB",x"22",x"EC",x"40",x"EB",x"CD",x"2C",x"1B", -- 0x1AB0
    x"C5",x"DC",x"E4",x"2B",x"D1",x"F1",x"D5",x"28", -- 0x1AB8
    x"27",x"D1",x"2A",x"F9",x"40",x"E3",x"C1",x"09", -- 0x1AC0
    x"E5",x"CD",x"55",x"19",x"E1",x"22",x"F9",x"40", -- 0x1AC8
    x"EB",x"74",x"D1",x"E5",x"23",x"23",x"73",x"23", -- 0x1AD0
    x"72",x"23",x"EB",x"2A",x"A7",x"40",x"EB",x"1B", -- 0x1AD8
    x"1B",x"1A",x"77",x"23",x"13",x"B7",x"20",x"F9", -- 0x1AE0
    x"D1",x"CD",x"FC",x"1A",x"CD",x"B5",x"41",x"CD", -- 0x1AE8
    x"5D",x"1B",x"CD",x"B8",x"41",x"C3",x"33",x"1A", -- 0x1AF0
    x"2A",x"A4",x"40",x"EB",x"62",x"6B",x"7E",x"23", -- 0x1AF8
    x"B6",x"C8",x"23",x"23",x"23",x"AF",x"BE",x"23", -- 0x1B00
    x"20",x"FC",x"EB",x"73",x"23",x"72",x"18",x"EC", -- 0x1B08
    x"11",x"00",x"00",x"D5",x"28",x"09",x"D1",x"CD", -- 0x1B10
    x"4F",x"1E",x"D5",x"28",x"0B",x"CF",x"CE",x"11", -- 0x1B18
    x"FA",x"FF",x"C4",x"4F",x"1E",x"C2",x"97",x"19", -- 0x1B20
    x"EB",x"D1",x"E3",x"E5",x"2A",x"A4",x"40",x"44", -- 0x1B28
    x"4D",x"7E",x"23",x"B6",x"2B",x"C8",x"23",x"23", -- 0x1B30
    x"7E",x"23",x"66",x"6F",x"DF",x"60",x"69",x"7E", -- 0x1B38
    x"23",x"66",x"6F",x"3F",x"C8",x"3F",x"D0",x"18", -- 0x1B40
    x"E6",x"C0",x"CD",x"C9",x"01",x"2A",x"A4",x"40", -- 0x1B48
    x"CD",x"F8",x"1D",x"32",x"E1",x"40",x"77",x"23", -- 0x1B50
    x"77",x"23",x"22",x"F9",x"40",x"2A",x"A4",x"40", -- 0x1B58
    x"2B",x"22",x"DF",x"40",x"06",x"1A",x"21",x"01", -- 0x1B60
    x"41",x"36",x"04",x"23",x"10",x"FB",x"AF",x"32", -- 0x1B68
    x"F2",x"40",x"6F",x"67",x"22",x"F0",x"40",x"22", -- 0x1B70
    x"F7",x"40",x"2A",x"B1",x"40",x"22",x"D6",x"40", -- 0x1B78
    x"CD",x"91",x"1D",x"2A",x"F9",x"40",x"22",x"FB", -- 0x1B80
    x"40",x"22",x"FD",x"40",x"CD",x"BB",x"41",x"C1", -- 0x1B88
    x"2A",x"A0",x"40",x"2B",x"2B",x"22",x"E8",x"40", -- 0x1B90
    x"23",x"23",x"F9",x"21",x"B5",x"40",x"22",x"B3", -- 0x1B98
    x"40",x"CD",x"8B",x"03",x"CD",x"69",x"21",x"AF", -- 0x1BA0
    x"67",x"6F",x"32",x"DC",x"40",x"E5",x"C5",x"2A", -- 0x1BA8
    x"DF",x"40",x"C9",x"3E",x"3F",x"CD",x"2A",x"03", -- 0x1BB0
    x"3E",x"20",x"CD",x"2A",x"03",x"C3",x"61",x"03", -- 0x1BB8
    x"AF",x"32",x"B0",x"40",x"4F",x"EB",x"2A",x"A7", -- 0x1BC0
    x"40",x"2B",x"2B",x"EB",x"7E",x"FE",x"20",x"CA", -- 0x1BC8
    x"5B",x"1C",x"47",x"FE",x"22",x"CA",x"77",x"1C", -- 0x1BD0
    x"B7",x"CA",x"7D",x"1C",x"3A",x"B0",x"40",x"B7", -- 0x1BD8
    x"7E",x"C2",x"5B",x"1C",x"FE",x"3F",x"3E",x"B2", -- 0x1BE0
    x"CA",x"5B",x"1C",x"7E",x"FE",x"30",x"38",x"05", -- 0x1BE8
    x"FE",x"3C",x"DA",x"5B",x"1C",x"D5",x"11",x"4F", -- 0x1BF0
    x"16",x"C5",x"01",x"3D",x"1C",x"C5",x"06",x"7F", -- 0x1BF8
    x"7E",x"FE",x"61",x"38",x"07",x"FE",x"7B",x"30", -- 0x1C00
    x"03",x"E6",x"5F",x"77",x"4E",x"EB",x"23",x"B6", -- 0x1C08
    x"F2",x"0E",x"1C",x"04",x"7E",x"CD",x"E2",x"38", -- 0x1C10
    x"B9",x"20",x"F3",x"EB",x"E5",x"13",x"1A",x"B7", -- 0x1C18
    x"FA",x"39",x"1C",x"4F",x"78",x"FE",x"8D",x"20", -- 0x1C20
    x"02",x"D7",x"2B",x"23",x"7E",x"FE",x"61",x"38", -- 0x1C28
    x"02",x"E6",x"5F",x"B9",x"28",x"E7",x"E1",x"18", -- 0x1C30
    x"D3",x"48",x"F1",x"EB",x"C9",x"EB",x"79",x"C1", -- 0x1C38
    x"D1",x"EB",x"FE",x"95",x"36",x"3A",x"20",x"02", -- 0x1C40
    x"0C",x"23",x"FE",x"FB",x"20",x"0C",x"36",x"3A", -- 0x1C48
    x"23",x"06",x"93",x"70",x"23",x"EB",x"0C",x"0C", -- 0x1C50
    x"18",x"1D",x"EB",x"23",x"12",x"13",x"0C",x"D6", -- 0x1C58
    x"3A",x"28",x"04",x"FE",x"4E",x"20",x"03",x"32", -- 0x1C60
    x"B0",x"40",x"D6",x"59",x"C2",x"CC",x"1B",x"47", -- 0x1C68
    x"7E",x"B7",x"28",x"09",x"B8",x"28",x"E4",x"23", -- 0x1C70
    x"12",x"0C",x"13",x"18",x"F3",x"21",x"05",x"00", -- 0x1C78
    x"44",x"09",x"44",x"4D",x"2A",x"A7",x"40",x"2B", -- 0x1C80
    x"2B",x"2B",x"12",x"13",x"12",x"13",x"12",x"C9", -- 0x1C88
    x"7C",x"92",x"C0",x"7D",x"93",x"C9",x"7E",x"E3", -- 0x1C90
    x"BE",x"23",x"E3",x"CA",x"78",x"1D",x"C3",x"97", -- 0x1C98
    x"19",x"3E",x"64",x"32",x"DC",x"40",x"CD",x"21", -- 0x1CA0
    x"1F",x"E3",x"CD",x"36",x"19",x"D1",x"20",x"05", -- 0x1CA8
    x"09",x"F9",x"22",x"E8",x"40",x"EB",x"0E",x"08", -- 0x1CB0
    x"CD",x"63",x"19",x"E5",x"CD",x"05",x"1F",x"E3", -- 0x1CB8
    x"E5",x"2A",x"A2",x"40",x"E3",x"CF",x"BD",x"E7", -- 0x1CC0
    x"CA",x"F6",x"0A",x"D2",x"F6",x"0A",x"F5",x"CD", -- 0x1CC8
    x"37",x"23",x"F1",x"E5",x"F2",x"EC",x"1C",x"CD", -- 0x1CD0
    x"7F",x"0A",x"E3",x"11",x"01",x"00",x"7E",x"FE", -- 0x1CD8
    x"CC",x"CC",x"01",x"2B",x"D5",x"E5",x"EB",x"CD", -- 0x1CE0
    x"9E",x"09",x"18",x"22",x"CD",x"B1",x"0A",x"CD", -- 0x1CE8
    x"BF",x"09",x"E1",x"C5",x"D5",x"01",x"00",x"81", -- 0x1CF0
    x"51",x"5A",x"7E",x"FE",x"CC",x"3E",x"01",x"20", -- 0x1CF8
    x"0E",x"CD",x"38",x"23",x"E5",x"CD",x"B1",x"0A", -- 0x1D00
    x"CD",x"BF",x"09",x"CD",x"55",x"09",x"E1",x"C5", -- 0x1D08
    x"D5",x"4F",x"E7",x"47",x"C5",x"E5",x"2A",x"DF", -- 0x1D10
    x"40",x"E3",x"06",x"81",x"C5",x"33",x"CD",x"58", -- 0x1D18
    x"03",x"B7",x"C4",x"A0",x"1D",x"22",x"E6",x"40", -- 0x1D20
    x"ED",x"73",x"E8",x"40",x"7E",x"FE",x"3A",x"28", -- 0x1D28
    x"29",x"B7",x"C2",x"97",x"19",x"23",x"7E",x"23", -- 0x1D30
    x"B6",x"CA",x"7E",x"19",x"23",x"5E",x"23",x"56", -- 0x1D38
    x"EB",x"22",x"A2",x"40",x"3A",x"1B",x"41",x"B7", -- 0x1D40
    x"28",x"0F",x"D5",x"3E",x"3C",x"CD",x"2A",x"03", -- 0x1D48
    x"CD",x"AF",x"0F",x"3E",x"3E",x"CD",x"2A",x"03", -- 0x1D50
    x"D1",x"EB",x"D7",x"11",x"1E",x"1D",x"D5",x"C8", -- 0x1D58
    x"D6",x"80",x"DA",x"21",x"1F",x"FE",x"3C",x"C3", -- 0x1D60
    x"C0",x"39",x"07",x"4F",x"06",x"00",x"EB",x"21", -- 0x1D68
    x"22",x"18",x"09",x"4E",x"23",x"46",x"C5",x"EB", -- 0x1D70
    x"23",x"7E",x"FE",x"3A",x"D0",x"FE",x"20",x"CA", -- 0x1D78
    x"78",x"1D",x"FE",x"0B",x"30",x"05",x"FE",x"09", -- 0x1D80
    x"D2",x"78",x"1D",x"FE",x"30",x"3F",x"3C",x"3D", -- 0x1D88
    x"C9",x"EB",x"2A",x"A4",x"40",x"2B",x"22",x"FF", -- 0x1D90
    x"40",x"EB",x"C9",x"CD",x"58",x"03",x"B7",x"C8", -- 0x1D98
    x"FE",x"60",x"CC",x"84",x"03",x"32",x"99",x"40", -- 0x1DA0
    x"3D",x"C0",x"3C",x"C3",x"B4",x"1D",x"C0",x"F5", -- 0x1DA8
    x"CC",x"BB",x"41",x"F1",x"22",x"E6",x"40",x"21", -- 0x1DB0
    x"B5",x"40",x"22",x"B3",x"40",x"21",x"F6",x"FF", -- 0x1DB8
    x"C1",x"2A",x"A2",x"40",x"E5",x"F5",x"7D",x"A4", -- 0x1DC0
    x"3C",x"28",x"09",x"22",x"F5",x"40",x"2A",x"E6", -- 0x1DC8
    x"40",x"22",x"F7",x"40",x"CD",x"8B",x"03",x"CD", -- 0x1DD0
    x"F9",x"20",x"F1",x"21",x"30",x"19",x"C2",x"06", -- 0x1DD8
    x"1A",x"C3",x"18",x"1A",x"2A",x"F7",x"40",x"7C", -- 0x1DE0
    x"B5",x"1E",x"20",x"CA",x"A2",x"19",x"EB",x"2A", -- 0x1DE8
    x"F5",x"40",x"CD",x"A0",x"38",x"EB",x"C9",x"3E", -- 0x1DF0
    x"AF",x"32",x"1B",x"41",x"C9",x"F1",x"E1",x"C9", -- 0x1DF8
    x"1E",x"03",x"01",x"1E",x"02",x"01",x"1E",x"04", -- 0x1E00
    x"01",x"1E",x"08",x"CD",x"3D",x"1E",x"01",x"97", -- 0x1E08
    x"19",x"C5",x"D8",x"D6",x"41",x"4F",x"47",x"D7", -- 0x1E10
    x"FE",x"CE",x"20",x"09",x"D7",x"CD",x"3D",x"1E", -- 0x1E18
    x"D8",x"D6",x"41",x"47",x"D7",x"78",x"91",x"D8", -- 0x1E20
    x"3C",x"E3",x"21",x"01",x"41",x"06",x"00",x"09", -- 0x1E28
    x"73",x"23",x"3D",x"20",x"FB",x"E1",x"7E",x"FE", -- 0x1E30
    x"2C",x"C0",x"D7",x"18",x"CE",x"7E",x"FE",x"41", -- 0x1E38
    x"D8",x"FE",x"5B",x"3F",x"C9",x"D7",x"CD",x"02", -- 0x1E40
    x"2B",x"F0",x"1E",x"08",x"C3",x"A2",x"19",x"7E", -- 0x1E48
    x"FE",x"2E",x"EB",x"2A",x"EC",x"40",x"EB",x"CA", -- 0x1E50
    x"78",x"1D",x"2B",x"11",x"00",x"00",x"D7",x"D0", -- 0x1E58
    x"E5",x"F5",x"21",x"98",x"19",x"DF",x"DA",x"97", -- 0x1E60
    x"19",x"62",x"6B",x"19",x"29",x"19",x"29",x"F1", -- 0x1E68
    x"D6",x"30",x"5F",x"16",x"00",x"19",x"EB",x"E1", -- 0x1E70
    x"18",x"E4",x"CA",x"61",x"1B",x"CD",x"46",x"1E", -- 0x1E78
    x"2B",x"D7",x"C0",x"E5",x"2A",x"B1",x"40",x"7D", -- 0x1E80
    x"93",x"5F",x"7C",x"9A",x"57",x"DA",x"7A",x"19", -- 0x1E88
    x"2A",x"F9",x"40",x"01",x"28",x"00",x"09",x"DF", -- 0x1E90
    x"D2",x"7A",x"19",x"EB",x"22",x"A0",x"40",x"E1", -- 0x1E98
    x"C3",x"61",x"1B",x"CA",x"5D",x"1B",x"CD",x"C7", -- 0x1EA0
    x"41",x"CD",x"61",x"1B",x"01",x"1E",x"1D",x"18", -- 0x1EA8
    x"10",x"0E",x"03",x"CD",x"63",x"19",x"C1",x"E5", -- 0x1EB0
    x"E5",x"2A",x"A2",x"40",x"E3",x"3E",x"91",x"F5", -- 0x1EB8
    x"33",x"C5",x"CD",x"5A",x"1E",x"CD",x"07",x"1F", -- 0x1EC0
    x"E5",x"2A",x"A2",x"40",x"DF",x"E1",x"23",x"DC", -- 0x1EC8
    x"2F",x"1B",x"D4",x"2C",x"1B",x"60",x"69",x"2B", -- 0x1ED0
    x"D8",x"1E",x"0E",x"C3",x"A2",x"19",x"C0",x"16", -- 0x1ED8
    x"FF",x"CD",x"36",x"19",x"F9",x"22",x"E8",x"40", -- 0x1EE0
    x"FE",x"91",x"1E",x"04",x"C2",x"A2",x"19",x"E1", -- 0x1EE8
    x"22",x"A2",x"40",x"23",x"7C",x"B5",x"20",x"07", -- 0x1EF0
    x"3A",x"DD",x"40",x"B7",x"C2",x"18",x"1A",x"21", -- 0x1EF8
    x"1E",x"1D",x"E3",x"3E",x"E1",x"01",x"3A",x"0E", -- 0x1F00
    x"00",x"06",x"00",x"79",x"48",x"47",x"7E",x"B7", -- 0x1F08
    x"C8",x"B8",x"C8",x"23",x"FE",x"22",x"28",x"F3", -- 0x1F10
    x"D6",x"8F",x"20",x"F2",x"B8",x"8A",x"57",x"18", -- 0x1F18
    x"ED",x"CD",x"0D",x"26",x"CF",x"D5",x"EB",x"22", -- 0x1F20
    x"DF",x"40",x"EB",x"D5",x"E7",x"F5",x"CD",x"37", -- 0x1F28
    x"23",x"F1",x"E3",x"C6",x"03",x"CD",x"19",x"28", -- 0x1F30
    x"CD",x"03",x"0A",x"E5",x"20",x"28",x"2A",x"21", -- 0x1F38
    x"41",x"E5",x"23",x"5E",x"23",x"56",x"2A",x"A4", -- 0x1F40
    x"40",x"DF",x"30",x"0E",x"2A",x"A0",x"40",x"DF", -- 0x1F48
    x"D1",x"30",x"0F",x"2A",x"F9",x"40",x"DF",x"30", -- 0x1F50
    x"09",x"3E",x"D1",x"CD",x"F5",x"29",x"EB",x"CD", -- 0x1F58
    x"43",x"28",x"CD",x"F5",x"29",x"E3",x"CD",x"D3", -- 0x1F60
    x"09",x"D1",x"E1",x"C9",x"FE",x"9E",x"20",x"25", -- 0x1F68
    x"D7",x"CF",x"8D",x"CD",x"5A",x"1E",x"7A",x"B3", -- 0x1F70
    x"28",x"09",x"CD",x"2A",x"1B",x"50",x"59",x"E1", -- 0x1F78
    x"D2",x"D9",x"1E",x"EB",x"22",x"F0",x"40",x"EB", -- 0x1F80
    x"D8",x"3A",x"F2",x"40",x"B7",x"C8",x"3A",x"9A", -- 0x1F88
    x"40",x"5F",x"C3",x"AB",x"19",x"CD",x"1C",x"2B", -- 0x1F90
    x"7E",x"47",x"FE",x"91",x"28",x"03",x"CF",x"8D", -- 0x1F98
    x"2B",x"4B",x"0D",x"78",x"CA",x"60",x"1D",x"CD", -- 0x1FA0
    x"5B",x"1E",x"FE",x"2C",x"C0",x"18",x"F3",x"11", -- 0x1FA8
    x"F2",x"40",x"1A",x"B7",x"CA",x"A0",x"19",x"3C", -- 0x1FB0
    x"32",x"9A",x"40",x"12",x"7E",x"FE",x"87",x"28", -- 0x1FB8
    x"0C",x"CD",x"5A",x"1E",x"C0",x"7A",x"B3",x"C2", -- 0x1FC0
    x"C5",x"1E",x"3C",x"18",x"02",x"D7",x"C0",x"2A", -- 0x1FC8
    x"EE",x"40",x"EB",x"2A",x"EA",x"40",x"22",x"A2", -- 0x1FD0
    x"40",x"EB",x"C0",x"7E",x"B7",x"20",x"04",x"23", -- 0x1FD8
    x"23",x"23",x"23",x"23",x"7A",x"A3",x"3C",x"C2", -- 0x1FE0
    x"05",x"1F",x"3A",x"DD",x"40",x"3D",x"CA",x"BE", -- 0x1FE8
    x"1D",x"C3",x"05",x"1F",x"CD",x"1C",x"2B",x"C0", -- 0x1FF0
    x"B7",x"CA",x"4A",x"1E",x"3D",x"87",x"5F",x"FE", -- 0x1FF8
    x"2D",x"38",x"02",x"1E",x"26",x"C3",x"A2",x"19", -- 0x2000
    x"11",x"0A",x"00",x"D5",x"28",x"17",x"CD",x"4F", -- 0x2008
    x"1E",x"EB",x"E3",x"28",x"11",x"EB",x"CF",x"2C", -- 0x2010
    x"EB",x"2A",x"E4",x"40",x"EB",x"28",x"06",x"CD", -- 0x2018
    x"5A",x"1E",x"C2",x"97",x"19",x"EB",x"7C",x"B5", -- 0x2020
    x"CA",x"4A",x"1E",x"22",x"E4",x"40",x"32",x"E1", -- 0x2028
    x"40",x"E1",x"22",x"E2",x"40",x"C1",x"C3",x"33", -- 0x2030
    x"1A",x"CD",x"37",x"23",x"7E",x"FE",x"2C",x"CC", -- 0x2038
    x"78",x"1D",x"FE",x"CA",x"CC",x"78",x"1D",x"2B", -- 0x2040
    x"E5",x"CD",x"94",x"09",x"E1",x"28",x"07",x"D7", -- 0x2048
    x"DA",x"C2",x"1E",x"C3",x"5F",x"1D",x"16",x"01", -- 0x2050
    x"CD",x"05",x"1F",x"B7",x"C8",x"D7",x"FE",x"95", -- 0x2058
    x"20",x"F6",x"15",x"20",x"F3",x"18",x"E8",x"3E", -- 0x2060
    x"01",x"32",x"9C",x"40",x"C3",x"9B",x"20",x"CD", -- 0x2068
    x"CA",x"41",x"FE",x"40",x"20",x"19",x"CD",x"01", -- 0x2070
    x"2B",x"E5",x"C3",x"D4",x"30",x"00",x"E5",x"21", -- 0x2078
    x"00",x"44",x"19",x"22",x"20",x"40",x"CD",x"2A", -- 0x2080
    x"36",x"32",x"A6",x"40",x"E1",x"CF",x"2C",x"FE", -- 0x2088
    x"23",x"20",x"08",x"CD",x"A9",x"35",x"3E",x"80", -- 0x2090
    x"32",x"9C",x"40",x"2B",x"D7",x"CC",x"FE",x"20", -- 0x2098
    x"CA",x"69",x"21",x"FE",x"BF",x"CA",x"BD",x"2C", -- 0x20A0
    x"FE",x"BC",x"CA",x"37",x"21",x"E5",x"FE",x"2C", -- 0x20A8
    x"CA",x"08",x"21",x"FE",x"3B",x"CA",x"64",x"21", -- 0x20B0
    x"C1",x"CD",x"37",x"23",x"E5",x"E7",x"28",x"32", -- 0x20B8
    x"CD",x"BD",x"0F",x"CD",x"65",x"28",x"CD",x"CD", -- 0x20C0
    x"41",x"2A",x"21",x"41",x"3A",x"9C",x"40",x"B7", -- 0x20C8
    x"FA",x"E9",x"20",x"28",x"08",x"3A",x"9B",x"40", -- 0x20D0
    x"86",x"FE",x"84",x"18",x"09",x"3A",x"9D",x"40", -- 0x20D8
    x"47",x"3A",x"A6",x"40",x"86",x"B8",x"D4",x"FE", -- 0x20E0
    x"20",x"CD",x"AA",x"28",x"3E",x"20",x"CD",x"2A", -- 0x20E8
    x"03",x"B7",x"CC",x"AA",x"28",x"E1",x"C3",x"9B", -- 0x20F0
    x"20",x"3A",x"A6",x"40",x"B7",x"C8",x"3E",x"0D", -- 0x20F8
    x"CD",x"2A",x"03",x"CD",x"D0",x"41",x"AF",x"C9", -- 0x2100
    x"CD",x"D3",x"41",x"3A",x"9C",x"40",x"B7",x"F2", -- 0x2108
    x"19",x"21",x"3E",x"2C",x"CD",x"2A",x"03",x"18", -- 0x2110
    x"4B",x"28",x"08",x"3A",x"9B",x"40",x"FE",x"70", -- 0x2118
    x"C3",x"2B",x"21",x"3A",x"9E",x"40",x"47",x"3A", -- 0x2120
    x"A6",x"40",x"B8",x"D4",x"FE",x"20",x"30",x"34", -- 0x2128
    x"D6",x"0A",x"30",x"FC",x"2F",x"18",x"23",x"CD", -- 0x2130
    x"1B",x"2B",x"CD",x"B2",x"30",x"CF",x"29",x"2B", -- 0x2138
    x"E5",x"CD",x"D3",x"41",x"3A",x"9C",x"40",x"B7", -- 0x2140
    x"FA",x"4A",x"1E",x"CA",x"53",x"21",x"3A",x"9B", -- 0x2148
    x"40",x"18",x"03",x"3A",x"A6",x"40",x"2F",x"83", -- 0x2150
    x"30",x"0A",x"3C",x"47",x"3E",x"20",x"CD",x"2A", -- 0x2158
    x"03",x"05",x"20",x"FA",x"E1",x"D7",x"C3",x"A0", -- 0x2160
    x"20",x"3A",x"9C",x"40",x"B7",x"00",x"00",x"00", -- 0x2168
    x"AF",x"32",x"9C",x"40",x"CD",x"BE",x"41",x"C9", -- 0x2170
    x"3F",x"52",x"45",x"44",x"4F",x"0D",x"00",x"3A", -- 0x2178
    x"DE",x"40",x"B7",x"C2",x"91",x"19",x"CD",x"B1", -- 0x2180
    x"30",x"B7",x"1E",x"2A",x"CA",x"A2",x"19",x"C1", -- 0x2188
    x"21",x"78",x"21",x"CD",x"A7",x"28",x"2A",x"E6", -- 0x2190
    x"40",x"C9",x"CD",x"28",x"28",x"7E",x"CD",x"D6", -- 0x2198
    x"41",x"D6",x"23",x"32",x"A9",x"40",x"7E",x"20", -- 0x21A0
    x"20",x"CD",x"AF",x"35",x"E5",x"06",x"FA",x"2A", -- 0x21A8
    x"A7",x"40",x"CD",x"ED",x"01",x"77",x"23",x"FE", -- 0x21B0
    x"0D",x"28",x"02",x"10",x"F5",x"2B",x"36",x"00", -- 0x21B8
    x"00",x"00",x"00",x"2A",x"A7",x"40",x"2B",x"18", -- 0x21C0
    x"22",x"01",x"DB",x"21",x"C5",x"FE",x"22",x"C0", -- 0x21C8
    x"CD",x"66",x"28",x"CF",x"3B",x"E5",x"CD",x"AA", -- 0x21D0
    x"28",x"E1",x"C9",x"E5",x"CD",x"B3",x"1B",x"C1", -- 0x21D8
    x"DA",x"BE",x"1D",x"23",x"7E",x"B7",x"2B",x"C5", -- 0x21E0
    x"CA",x"04",x"1F",x"36",x"2C",x"18",x"05",x"E5", -- 0x21E8
    x"2A",x"FF",x"40",x"F6",x"AF",x"32",x"DE",x"40", -- 0x21F0
    x"E3",x"18",x"02",x"CF",x"2C",x"CD",x"0D",x"26", -- 0x21F8
    x"E3",x"D5",x"7E",x"FE",x"2C",x"28",x"26",x"3A", -- 0x2200
    x"DE",x"40",x"B7",x"C2",x"96",x"22",x"3A",x"A9", -- 0x2208
    x"40",x"B7",x"1E",x"06",x"CA",x"A2",x"19",x"3E", -- 0x2210
    x"3F",x"CD",x"2A",x"03",x"CD",x"B3",x"1B",x"D1", -- 0x2218
    x"C1",x"DA",x"BE",x"1D",x"23",x"7E",x"B7",x"2B", -- 0x2220
    x"C5",x"CA",x"04",x"1F",x"D5",x"CD",x"DC",x"41", -- 0x2228
    x"E7",x"F5",x"20",x"19",x"D7",x"57",x"47",x"FE", -- 0x2230
    x"22",x"28",x"05",x"16",x"3A",x"06",x"2C",x"2B", -- 0x2238
    x"CD",x"69",x"28",x"F1",x"EB",x"21",x"5A",x"22", -- 0x2240
    x"E3",x"D5",x"C3",x"33",x"1F",x"D7",x"F1",x"F5", -- 0x2248
    x"01",x"43",x"22",x"C5",x"DA",x"6C",x"0E",x"D2", -- 0x2250
    x"65",x"0E",x"2B",x"D7",x"28",x"05",x"FE",x"2C", -- 0x2258
    x"C2",x"7F",x"21",x"E3",x"2B",x"D7",x"C2",x"FB", -- 0x2260
    x"21",x"D1",x"00",x"00",x"00",x"00",x"00",x"3A", -- 0x2268
    x"DE",x"40",x"B7",x"EB",x"C2",x"96",x"1D",x"D5", -- 0x2270
    x"CD",x"DF",x"41",x"B6",x"21",x"86",x"22",x"C4", -- 0x2278
    x"A7",x"28",x"E1",x"C3",x"69",x"21",x"3F",x"45", -- 0x2280
    x"78",x"74",x"72",x"61",x"20",x"69",x"67",x"6E", -- 0x2288
    x"6F",x"72",x"65",x"64",x"0D",x"00",x"CD",x"05", -- 0x2290
    x"1F",x"B7",x"20",x"12",x"23",x"7E",x"23",x"B6", -- 0x2298
    x"1E",x"06",x"CA",x"A2",x"19",x"23",x"5E",x"23", -- 0x22A0
    x"56",x"EB",x"22",x"DA",x"40",x"EB",x"D7",x"FE", -- 0x22A8
    x"88",x"20",x"E3",x"C3",x"2D",x"22",x"11",x"00", -- 0x22B0
    x"00",x"C4",x"0D",x"26",x"22",x"DF",x"40",x"CD", -- 0x22B8
    x"36",x"19",x"C2",x"9D",x"19",x"F9",x"22",x"E8", -- 0x22C0
    x"40",x"D5",x"7E",x"23",x"F5",x"D5",x"7E",x"23", -- 0x22C8
    x"B7",x"FA",x"EA",x"22",x"CD",x"B1",x"09",x"E3", -- 0x22D0
    x"E5",x"CD",x"0B",x"07",x"E1",x"CD",x"CB",x"09", -- 0x22D8
    x"E1",x"CD",x"C2",x"09",x"E5",x"CD",x"0C",x"0A", -- 0x22E0
    x"18",x"29",x"23",x"23",x"23",x"23",x"4E",x"23", -- 0x22E8
    x"46",x"23",x"E3",x"5E",x"23",x"56",x"E5",x"69", -- 0x22F0
    x"60",x"CD",x"D2",x"0B",x"3A",x"AF",x"40",x"FE", -- 0x22F8
    x"04",x"CA",x"B2",x"07",x"EB",x"E1",x"72",x"2B", -- 0x2300
    x"73",x"E1",x"D5",x"5E",x"23",x"56",x"23",x"E3", -- 0x2308
    x"CD",x"39",x"0A",x"E1",x"C1",x"90",x"CD",x"C2", -- 0x2310
    x"09",x"28",x"09",x"EB",x"22",x"A2",x"40",x"69", -- 0x2318
    x"60",x"C3",x"1A",x"1D",x"F9",x"22",x"E8",x"40", -- 0x2320
    x"2A",x"DF",x"40",x"7E",x"FE",x"2C",x"C2",x"1E", -- 0x2328
    x"1D",x"D7",x"CD",x"B9",x"22",x"CF",x"28",x"2B", -- 0x2330
    x"16",x"00",x"D5",x"0E",x"01",x"CD",x"63",x"19", -- 0x2338
    x"CD",x"9F",x"24",x"22",x"F3",x"40",x"2A",x"F3", -- 0x2340
    x"40",x"C1",x"7E",x"16",x"00",x"D6",x"D4",x"38", -- 0x2348
    x"13",x"FE",x"03",x"30",x"0F",x"FE",x"01",x"17", -- 0x2350
    x"AA",x"BA",x"57",x"DA",x"97",x"19",x"22",x"D8", -- 0x2358
    x"40",x"D7",x"18",x"E9",x"7A",x"B7",x"C2",x"EC", -- 0x2360
    x"23",x"7E",x"22",x"D8",x"40",x"D6",x"CD",x"D8", -- 0x2368
    x"FE",x"07",x"D0",x"5F",x"3A",x"AF",x"40",x"D6", -- 0x2370
    x"03",x"B3",x"CA",x"8F",x"29",x"21",x"9A",x"18", -- 0x2378
    x"19",x"78",x"56",x"BA",x"D0",x"C5",x"01",x"46", -- 0x2380
    x"23",x"C5",x"7A",x"FE",x"7F",x"CA",x"D4",x"23", -- 0x2388
    x"FE",x"51",x"DA",x"E1",x"23",x"21",x"21",x"41", -- 0x2390
    x"B7",x"3A",x"AF",x"40",x"3D",x"3D",x"3D",x"CA", -- 0x2398
    x"F6",x"0A",x"4E",x"23",x"46",x"C5",x"FA",x"C5", -- 0x23A0
    x"23",x"23",x"4E",x"23",x"46",x"C5",x"F5",x"B7", -- 0x23A8
    x"E2",x"C4",x"23",x"F1",x"23",x"38",x"03",x"21", -- 0x23B0
    x"1D",x"41",x"4E",x"23",x"46",x"23",x"C5",x"4E", -- 0x23B8
    x"23",x"46",x"C5",x"06",x"F1",x"C6",x"03",x"4B", -- 0x23C0
    x"47",x"C5",x"01",x"06",x"24",x"C5",x"2A",x"D8", -- 0x23C8
    x"40",x"C3",x"3A",x"23",x"CD",x"B1",x"0A",x"CD", -- 0x23D0
    x"A4",x"09",x"01",x"F2",x"13",x"16",x"7F",x"18", -- 0x23D8
    x"EC",x"D5",x"CD",x"7F",x"0A",x"D1",x"E5",x"01", -- 0x23E0
    x"E9",x"25",x"18",x"E1",x"78",x"FE",x"64",x"D0", -- 0x23E8
    x"C5",x"D5",x"11",x"04",x"64",x"21",x"B8",x"25", -- 0x23F0
    x"E5",x"E7",x"C2",x"95",x"23",x"2A",x"21",x"41", -- 0x23F8
    x"E5",x"01",x"8C",x"25",x"18",x"C7",x"C1",x"79", -- 0x2400
    x"32",x"B0",x"40",x"78",x"FE",x"08",x"28",x"28", -- 0x2408
    x"3A",x"AF",x"40",x"FE",x"08",x"CA",x"60",x"24", -- 0x2410
    x"57",x"78",x"FE",x"04",x"CA",x"72",x"24",x"7A", -- 0x2418
    x"FE",x"03",x"CA",x"F6",x"0A",x"D2",x"7C",x"24", -- 0x2420
    x"21",x"BF",x"18",x"06",x"00",x"09",x"09",x"4E", -- 0x2428
    x"23",x"46",x"D1",x"2A",x"21",x"41",x"C5",x"C9", -- 0x2430
    x"CD",x"DB",x"0A",x"CD",x"FC",x"09",x"E1",x"22", -- 0x2438
    x"1F",x"41",x"E1",x"22",x"1D",x"41",x"C1",x"D1", -- 0x2440
    x"CD",x"B4",x"09",x"CD",x"DB",x"0A",x"21",x"AB", -- 0x2448
    x"18",x"3A",x"B0",x"40",x"07",x"C5",x"4F",x"06", -- 0x2450
    x"00",x"09",x"C1",x"7E",x"23",x"66",x"6F",x"E9", -- 0x2458
    x"C5",x"CD",x"FC",x"09",x"F1",x"32",x"AF",x"40", -- 0x2460
    x"FE",x"04",x"28",x"DA",x"E1",x"22",x"21",x"41", -- 0x2468
    x"18",x"D9",x"CD",x"B1",x"0A",x"C1",x"D1",x"21", -- 0x2470
    x"B5",x"18",x"18",x"D5",x"E1",x"CD",x"A4",x"09", -- 0x2478
    x"CD",x"CF",x"0A",x"CD",x"BF",x"09",x"E1",x"22", -- 0x2480
    x"23",x"41",x"E1",x"22",x"21",x"41",x"18",x"E7", -- 0x2488
    x"E5",x"EB",x"CD",x"CF",x"0A",x"E1",x"CD",x"A4", -- 0x2490
    x"09",x"CD",x"CF",x"0A",x"C3",x"A0",x"08",x"D7", -- 0x2498
    x"1E",x"28",x"CA",x"A2",x"19",x"DA",x"6C",x"0E", -- 0x24A0
    x"CD",x"3D",x"1E",x"D2",x"40",x"25",x"FE",x"CD", -- 0x24A8
    x"28",x"ED",x"FE",x"2E",x"CA",x"6C",x"0E",x"FE", -- 0x24B0
    x"CE",x"CA",x"32",x"25",x"FE",x"22",x"CA",x"66", -- 0x24B8
    x"28",x"FE",x"CB",x"CA",x"C4",x"25",x"FE",x"26", -- 0x24C0
    x"CA",x"E3",x"34",x"FE",x"C3",x"20",x"0A",x"D7", -- 0x24C8
    x"3A",x"9A",x"40",x"E5",x"CD",x"F8",x"27",x"E1", -- 0x24D0
    x"C9",x"FE",x"C2",x"20",x"0A",x"D7",x"E5",x"2A", -- 0x24D8
    x"EA",x"40",x"CD",x"66",x"0C",x"E1",x"C9",x"FE", -- 0x24E0
    x"C0",x"20",x"14",x"D7",x"CF",x"28",x"CD",x"0D", -- 0x24E8
    x"26",x"CF",x"29",x"E5",x"EB",x"7C",x"B5",x"CA", -- 0x24F0
    x"4A",x"1E",x"CD",x"9A",x"0A",x"E1",x"C9",x"FE", -- 0x24F8
    x"C1",x"C3",x"7A",x"3F",x"FE",x"C5",x"CA",x"9D", -- 0x2500
    x"41",x"FE",x"C8",x"CA",x"C9",x"27",x"FE",x"C7", -- 0x2508
    x"CA",x"76",x"41",x"FE",x"C6",x"CA",x"32",x"01", -- 0x2510
    x"FE",x"C9",x"CA",x"9D",x"01",x"FE",x"C4",x"CA", -- 0x2518
    x"2F",x"2A",x"FE",x"BE",x"CA",x"55",x"41",x"D6", -- 0x2520
    x"D7",x"D2",x"4E",x"25",x"CD",x"35",x"23",x"CF", -- 0x2528
    x"29",x"C9",x"16",x"7D",x"CD",x"3A",x"23",x"2A", -- 0x2530
    x"F3",x"40",x"E5",x"CD",x"7B",x"09",x"E1",x"C9", -- 0x2538
    x"CD",x"0D",x"26",x"E5",x"EB",x"22",x"21",x"41", -- 0x2540
    x"E7",x"C4",x"F7",x"09",x"E1",x"C9",x"06",x"00", -- 0x2548
    x"07",x"4F",x"C5",x"D7",x"79",x"FE",x"41",x"38", -- 0x2550
    x"16",x"CD",x"35",x"23",x"CF",x"2C",x"CD",x"F4", -- 0x2558
    x"0A",x"EB",x"2A",x"21",x"41",x"E3",x"E5",x"EB", -- 0x2560
    x"CD",x"1C",x"2B",x"EB",x"E3",x"18",x"14",x"CD", -- 0x2568
    x"2C",x"25",x"E3",x"7D",x"FE",x"0C",x"38",x"07", -- 0x2570
    x"FE",x"1B",x"E5",x"DC",x"B1",x"0A",x"E1",x"11", -- 0x2578
    x"3E",x"25",x"D5",x"01",x"08",x"16",x"09",x"4E", -- 0x2580
    x"23",x"66",x"69",x"E9",x"CD",x"D7",x"29",x"7E", -- 0x2588
    x"23",x"4E",x"23",x"46",x"D1",x"C5",x"F5",x"CD", -- 0x2590
    x"DE",x"29",x"D1",x"5E",x"23",x"4E",x"23",x"46", -- 0x2598
    x"E1",x"7B",x"B2",x"C8",x"7A",x"D6",x"01",x"D8", -- 0x25A0
    x"AF",x"BB",x"3C",x"D0",x"15",x"1D",x"0A",x"BE", -- 0x25A8
    x"23",x"03",x"28",x"ED",x"3F",x"C3",x"60",x"09", -- 0x25B0
    x"3C",x"8F",x"C1",x"A0",x"C6",x"FF",x"9F",x"CD", -- 0x25B8
    x"8D",x"09",x"18",x"12",x"16",x"5A",x"CD",x"3A", -- 0x25C0
    x"23",x"CD",x"7F",x"0A",x"7D",x"2F",x"6F",x"7C", -- 0x25C8
    x"2F",x"67",x"22",x"21",x"41",x"C1",x"C3",x"46", -- 0x25D0
    x"23",x"3A",x"AF",x"40",x"FE",x"08",x"30",x"05", -- 0x25D8
    x"D6",x"03",x"B7",x"37",x"C9",x"D6",x"03",x"B7", -- 0x25E0
    x"C9",x"C5",x"CD",x"7F",x"0A",x"F1",x"D1",x"01", -- 0x25E8
    x"FA",x"27",x"C5",x"FE",x"46",x"20",x"06",x"7B", -- 0x25F0
    x"B5",x"6F",x"7C",x"B2",x"C9",x"7B",x"A5",x"6F", -- 0x25F8
    x"7C",x"A2",x"C9",x"2B",x"D7",x"C8",x"CF",x"2C", -- 0x2600
    x"01",x"03",x"26",x"C5",x"F6",x"AF",x"32",x"AE", -- 0x2608
    x"40",x"46",x"CD",x"3D",x"1E",x"DA",x"97",x"19", -- 0x2610
    x"AF",x"4F",x"D7",x"38",x"05",x"CD",x"3D",x"1E", -- 0x2618
    x"38",x"09",x"4F",x"D7",x"38",x"FD",x"CD",x"3D", -- 0x2620
    x"1E",x"30",x"F8",x"11",x"52",x"26",x"D5",x"16", -- 0x2628
    x"02",x"FE",x"25",x"C8",x"14",x"FE",x"24",x"C8", -- 0x2630
    x"14",x"FE",x"21",x"C8",x"16",x"08",x"FE",x"23", -- 0x2638
    x"C8",x"78",x"D6",x"41",x"E6",x"7F",x"5F",x"16", -- 0x2640
    x"00",x"E5",x"21",x"01",x"41",x"19",x"56",x"E1", -- 0x2648
    x"2B",x"C9",x"7A",x"32",x"AF",x"40",x"D7",x"3A", -- 0x2650
    x"DC",x"40",x"B7",x"C2",x"64",x"26",x"7E",x"D6", -- 0x2658
    x"28",x"CA",x"E9",x"26",x"AF",x"32",x"DC",x"40", -- 0x2660
    x"E5",x"D5",x"2A",x"F9",x"40",x"EB",x"2A",x"FB", -- 0x2668
    x"40",x"DF",x"E1",x"28",x"19",x"1A",x"6F",x"BC", -- 0x2670
    x"13",x"20",x"0B",x"1A",x"B9",x"20",x"07",x"13", -- 0x2678
    x"1A",x"B8",x"CA",x"CC",x"26",x"3E",x"13",x"13", -- 0x2680
    x"E5",x"26",x"00",x"19",x"18",x"DF",x"7C",x"E1", -- 0x2688
    x"E3",x"F5",x"D5",x"11",x"F1",x"24",x"DF",x"28", -- 0x2690
    x"36",x"11",x"43",x"25",x"DF",x"D1",x"28",x"35", -- 0x2698
    x"F1",x"E3",x"E5",x"C5",x"4F",x"06",x"00",x"C5", -- 0x26A0
    x"03",x"03",x"03",x"2A",x"FD",x"40",x"E5",x"09", -- 0x26A8
    x"C1",x"E5",x"CD",x"55",x"19",x"E1",x"22",x"FD", -- 0x26B0
    x"40",x"60",x"69",x"22",x"FB",x"40",x"2B",x"36", -- 0x26B8
    x"00",x"DF",x"20",x"FA",x"D1",x"73",x"23",x"D1", -- 0x26C0
    x"73",x"23",x"72",x"EB",x"13",x"E1",x"C9",x"57", -- 0x26C8
    x"5F",x"F1",x"F1",x"E3",x"C9",x"32",x"24",x"41", -- 0x26D0
    x"C1",x"67",x"6F",x"22",x"21",x"41",x"E7",x"20", -- 0x26D8
    x"06",x"21",x"28",x"19",x"22",x"21",x"41",x"E1", -- 0x26E0
    x"C9",x"E5",x"2A",x"AE",x"40",x"E3",x"57",x"D5", -- 0x26E8
    x"C5",x"CD",x"45",x"1E",x"C1",x"F1",x"EB",x"E3", -- 0x26F0
    x"E5",x"EB",x"3C",x"57",x"7E",x"FE",x"2C",x"28", -- 0x26F8
    x"EE",x"CF",x"29",x"22",x"F3",x"40",x"E1",x"22", -- 0x2700
    x"AE",x"40",x"D5",x"2A",x"FB",x"40",x"3E",x"19", -- 0x2708
    x"EB",x"2A",x"FD",x"40",x"EB",x"DF",x"3A",x"AF", -- 0x2710
    x"40",x"28",x"27",x"BE",x"23",x"20",x"08",x"7E", -- 0x2718
    x"B9",x"23",x"20",x"04",x"7E",x"B8",x"3E",x"23", -- 0x2720
    x"23",x"5E",x"23",x"56",x"23",x"20",x"E0",x"3A", -- 0x2728
    x"AE",x"40",x"B7",x"1E",x"12",x"C2",x"A2",x"19", -- 0x2730
    x"F1",x"96",x"CA",x"95",x"27",x"1E",x"10",x"C3", -- 0x2738
    x"A2",x"19",x"77",x"23",x"5F",x"16",x"00",x"F1", -- 0x2740
    x"71",x"23",x"70",x"23",x"4F",x"CD",x"63",x"19", -- 0x2748
    x"23",x"23",x"22",x"D8",x"40",x"71",x"23",x"3A", -- 0x2750
    x"AE",x"40",x"17",x"79",x"01",x"0B",x"00",x"30", -- 0x2758
    x"02",x"C1",x"03",x"71",x"23",x"70",x"23",x"F5", -- 0x2760
    x"CD",x"AA",x"0B",x"F1",x"3D",x"20",x"ED",x"F5", -- 0x2768
    x"42",x"4B",x"EB",x"19",x"38",x"C7",x"CD",x"6C", -- 0x2770
    x"19",x"22",x"FD",x"40",x"2B",x"36",x"00",x"DF", -- 0x2778
    x"20",x"FA",x"03",x"57",x"2A",x"D8",x"40",x"5E", -- 0x2780
    x"EB",x"29",x"09",x"EB",x"2B",x"2B",x"73",x"23", -- 0x2788
    x"72",x"23",x"F1",x"38",x"30",x"47",x"4F",x"7E", -- 0x2790
    x"23",x"16",x"E1",x"5E",x"23",x"56",x"23",x"E3", -- 0x2798
    x"F5",x"DF",x"D2",x"3D",x"27",x"CD",x"AA",x"0B", -- 0x27A0
    x"19",x"F1",x"3D",x"44",x"4D",x"20",x"EB",x"3A", -- 0x27A8
    x"AF",x"40",x"44",x"4D",x"29",x"D6",x"04",x"38", -- 0x27B0
    x"04",x"29",x"28",x"06",x"29",x"B7",x"E2",x"C2", -- 0x27B8
    x"27",x"09",x"C1",x"09",x"EB",x"2A",x"F3",x"40", -- 0x27C0
    x"C9",x"AF",x"E5",x"32",x"AF",x"40",x"CD",x"D4", -- 0x27C8
    x"27",x"E1",x"D7",x"C9",x"2A",x"FD",x"40",x"EB", -- 0x27D0
    x"21",x"00",x"00",x"39",x"E7",x"20",x"0D",x"CD", -- 0x27D8
    x"DA",x"29",x"CD",x"E6",x"28",x"2A",x"A0",x"40", -- 0x27E0
    x"EB",x"2A",x"D6",x"40",x"7D",x"93",x"6F",x"7C", -- 0x27E8
    x"9A",x"67",x"C3",x"66",x"0C",x"3A",x"A6",x"40", -- 0x27F0
    x"6F",x"AF",x"67",x"C3",x"9A",x"0A",x"CD",x"A9", -- 0x27F8
    x"41",x"D7",x"CD",x"2C",x"25",x"E5",x"21",x"90", -- 0x2800
    x"08",x"E5",x"3A",x"AF",x"40",x"F5",x"FE",x"03", -- 0x2808
    x"CC",x"DA",x"29",x"F1",x"EB",x"2A",x"8E",x"40", -- 0x2810
    x"E9",x"E5",x"E6",x"07",x"21",x"A1",x"18",x"4F", -- 0x2818
    x"06",x"00",x"09",x"CD",x"86",x"25",x"E1",x"C9", -- 0x2820
    x"E5",x"2A",x"A2",x"40",x"23",x"7C",x"B5",x"E1", -- 0x2828
    x"C0",x"1E",x"16",x"C3",x"A2",x"19",x"CD",x"BD", -- 0x2830
    x"0F",x"CD",x"65",x"28",x"CD",x"DA",x"29",x"01", -- 0x2838
    x"2B",x"2A",x"C5",x"7E",x"23",x"E5",x"CD",x"BF", -- 0x2840
    x"28",x"E1",x"4E",x"23",x"46",x"CD",x"5A",x"28", -- 0x2848
    x"E5",x"6F",x"CD",x"CE",x"29",x"D1",x"C9",x"CD", -- 0x2850
    x"BF",x"28",x"21",x"D3",x"40",x"E5",x"77",x"23", -- 0x2858
    x"73",x"23",x"72",x"E1",x"C9",x"2B",x"06",x"22", -- 0x2860
    x"50",x"E5",x"0E",x"FF",x"23",x"7E",x"0C",x"B7", -- 0x2868
    x"28",x"06",x"BA",x"28",x"03",x"B8",x"20",x"F4", -- 0x2870
    x"FE",x"22",x"CC",x"78",x"1D",x"E3",x"23",x"EB", -- 0x2878
    x"79",x"CD",x"5A",x"28",x"11",x"D3",x"40",x"3E", -- 0x2880
    x"D5",x"2A",x"B3",x"40",x"22",x"21",x"41",x"3E", -- 0x2888
    x"03",x"32",x"AF",x"40",x"CD",x"D3",x"09",x"11", -- 0x2890
    x"D6",x"40",x"DF",x"22",x"B3",x"40",x"E1",x"7E", -- 0x2898
    x"C0",x"1E",x"1E",x"C3",x"A2",x"19",x"23",x"CD", -- 0x28A0
    x"65",x"28",x"CD",x"DA",x"29",x"CD",x"C4",x"09", -- 0x28A8
    x"14",x"15",x"C8",x"0A",x"CD",x"2A",x"03",x"FE", -- 0x28B0
    x"0D",x"CC",x"03",x"21",x"03",x"18",x"F2",x"B7", -- 0x28B8
    x"0E",x"F1",x"F5",x"2A",x"A0",x"40",x"EB",x"2A", -- 0x28C0
    x"D6",x"40",x"2F",x"4F",x"06",x"FF",x"09",x"23", -- 0x28C8
    x"DF",x"38",x"07",x"22",x"D6",x"40",x"23",x"EB", -- 0x28D0
    x"F1",x"C9",x"F1",x"1E",x"1A",x"CA",x"A2",x"19", -- 0x28D8
    x"BF",x"F5",x"01",x"C1",x"28",x"C5",x"2A",x"B1", -- 0x28E0
    x"40",x"22",x"D6",x"40",x"21",x"00",x"00",x"E5", -- 0x28E8
    x"2A",x"A0",x"40",x"E5",x"21",x"B5",x"40",x"EB", -- 0x28F0
    x"2A",x"B3",x"40",x"EB",x"DF",x"01",x"F7",x"28", -- 0x28F8
    x"C2",x"4A",x"29",x"2A",x"F9",x"40",x"EB",x"2A", -- 0x2900
    x"FB",x"40",x"EB",x"DF",x"28",x"13",x"7E",x"23", -- 0x2908
    x"23",x"23",x"FE",x"03",x"20",x"04",x"CD",x"4B", -- 0x2910
    x"29",x"AF",x"5F",x"16",x"00",x"19",x"18",x"E6", -- 0x2918
    x"C1",x"EB",x"2A",x"FD",x"40",x"EB",x"DF",x"CA", -- 0x2920
    x"6B",x"29",x"7E",x"23",x"CD",x"C2",x"09",x"E5", -- 0x2928
    x"09",x"FE",x"03",x"20",x"EB",x"22",x"D8",x"40", -- 0x2930
    x"E1",x"4E",x"06",x"00",x"09",x"09",x"23",x"EB", -- 0x2938
    x"2A",x"D8",x"40",x"EB",x"DF",x"28",x"DA",x"01", -- 0x2940
    x"3F",x"29",x"C5",x"AF",x"B6",x"23",x"5E",x"23", -- 0x2948
    x"56",x"23",x"C8",x"44",x"4D",x"2A",x"D6",x"40", -- 0x2950
    x"DF",x"60",x"69",x"D8",x"E1",x"E3",x"DF",x"E3", -- 0x2958
    x"E5",x"60",x"69",x"D0",x"C1",x"F1",x"F1",x"E5", -- 0x2960
    x"D5",x"C5",x"C9",x"D1",x"E1",x"7D",x"B4",x"C8", -- 0x2968
    x"2B",x"46",x"2B",x"4E",x"E5",x"2B",x"6E",x"26", -- 0x2970
    x"00",x"09",x"50",x"59",x"2B",x"44",x"4D",x"2A", -- 0x2978
    x"D6",x"40",x"CD",x"58",x"19",x"E1",x"71",x"23", -- 0x2980
    x"70",x"69",x"60",x"2B",x"C3",x"E9",x"28",x"C5", -- 0x2988
    x"E5",x"2A",x"21",x"41",x"E3",x"CD",x"9F",x"24", -- 0x2990
    x"E3",x"CD",x"F4",x"0A",x"7E",x"E5",x"2A",x"21", -- 0x2998
    x"41",x"E5",x"86",x"1E",x"1C",x"DA",x"A2",x"19", -- 0x29A0
    x"CD",x"57",x"28",x"D1",x"CD",x"DE",x"29",x"E3", -- 0x29A8
    x"CD",x"DD",x"29",x"E5",x"2A",x"D4",x"40",x"EB", -- 0x29B0
    x"CD",x"C6",x"29",x"CD",x"C6",x"29",x"21",x"49", -- 0x29B8
    x"23",x"E3",x"E5",x"C3",x"84",x"28",x"E1",x"E3", -- 0x29C0
    x"7E",x"23",x"4E",x"23",x"46",x"6F",x"2C",x"2D", -- 0x29C8
    x"C8",x"0A",x"12",x"03",x"13",x"18",x"F8",x"CD", -- 0x29D0
    x"F4",x"0A",x"2A",x"21",x"41",x"EB",x"CD",x"F5", -- 0x29D8
    x"29",x"EB",x"C0",x"D5",x"50",x"59",x"1B",x"4E", -- 0x29E0
    x"2A",x"D6",x"40",x"DF",x"20",x"05",x"47",x"09", -- 0x29E8
    x"22",x"D6",x"40",x"E1",x"C9",x"2A",x"B3",x"40", -- 0x29F0
    x"2B",x"46",x"2B",x"4E",x"2B",x"DF",x"C0",x"22", -- 0x29F8
    x"B3",x"40",x"C9",x"01",x"F8",x"27",x"C5",x"CD", -- 0x2A00
    x"D7",x"29",x"AF",x"57",x"7E",x"B7",x"C9",x"01", -- 0x2A08
    x"F8",x"27",x"C5",x"CD",x"07",x"2A",x"CA",x"4A", -- 0x2A10
    x"1E",x"23",x"5E",x"23",x"56",x"1A",x"C9",x"3E", -- 0x2A18
    x"01",x"CD",x"57",x"28",x"CD",x"1F",x"2B",x"2A", -- 0x2A20
    x"D4",x"40",x"73",x"C1",x"C3",x"84",x"28",x"D7", -- 0x2A28
    x"CF",x"28",x"CD",x"1C",x"2B",x"D5",x"CF",x"2C", -- 0x2A30
    x"CD",x"37",x"23",x"CF",x"29",x"E3",x"E5",x"E7", -- 0x2A38
    x"28",x"05",x"CD",x"1F",x"2B",x"18",x"03",x"CD", -- 0x2A40
    x"13",x"2A",x"D1",x"F5",x"F5",x"7B",x"CD",x"57", -- 0x2A48
    x"28",x"5F",x"F1",x"1C",x"1D",x"28",x"D4",x"2A", -- 0x2A50
    x"D4",x"40",x"77",x"23",x"1D",x"20",x"FB",x"18", -- 0x2A58
    x"CA",x"CD",x"DF",x"2A",x"AF",x"E3",x"4F",x"3E", -- 0x2A60
    x"E5",x"E5",x"7E",x"B8",x"38",x"02",x"78",x"11", -- 0x2A68
    x"0E",x"00",x"C5",x"CD",x"BF",x"28",x"C1",x"E1", -- 0x2A70
    x"E5",x"23",x"46",x"23",x"66",x"68",x"06",x"00", -- 0x2A78
    x"09",x"44",x"4D",x"CD",x"5A",x"28",x"6F",x"CD", -- 0x2A80
    x"CE",x"29",x"D1",x"CD",x"DE",x"29",x"C3",x"84", -- 0x2A88
    x"28",x"CD",x"DF",x"2A",x"D1",x"D5",x"1A",x"90", -- 0x2A90
    x"18",x"CB",x"EB",x"7E",x"CD",x"E2",x"2A",x"04", -- 0x2A98
    x"05",x"CA",x"4A",x"1E",x"C5",x"1E",x"FF",x"FE", -- 0x2AA0
    x"29",x"28",x"05",x"CF",x"2C",x"CD",x"1C",x"2B", -- 0x2AA8
    x"CF",x"29",x"F1",x"E3",x"01",x"69",x"2A",x"C5", -- 0x2AB0
    x"3D",x"BE",x"06",x"00",x"D0",x"4F",x"7E",x"91", -- 0x2AB8
    x"BB",x"47",x"D8",x"43",x"C9",x"CD",x"07",x"2A", -- 0x2AC0
    x"CA",x"F8",x"27",x"5F",x"23",x"7E",x"23",x"66", -- 0x2AC8
    x"6F",x"E5",x"19",x"46",x"72",x"E3",x"C5",x"7E", -- 0x2AD0
    x"CD",x"65",x"0E",x"C1",x"E1",x"70",x"C9",x"EB", -- 0x2AD8
    x"CF",x"29",x"C1",x"D1",x"C5",x"43",x"C9",x"FE", -- 0x2AE0
    x"7A",x"C2",x"97",x"19",x"C3",x"D9",x"41",x"CD", -- 0x2AE8
    x"1F",x"2B",x"32",x"94",x"40",x"CD",x"93",x"40", -- 0x2AF0
    x"C3",x"F8",x"27",x"CD",x"0E",x"2B",x"C3",x"96", -- 0x2AF8
    x"40",x"D7",x"CD",x"37",x"23",x"E5",x"CD",x"7F", -- 0x2B00
    x"0A",x"EB",x"E1",x"7A",x"B7",x"C9",x"CD",x"1C", -- 0x2B08
    x"2B",x"32",x"94",x"40",x"32",x"97",x"40",x"CF", -- 0x2B10
    x"2C",x"18",x"01",x"D7",x"CD",x"37",x"23",x"CD", -- 0x2B18
    x"05",x"2B",x"C2",x"4A",x"1E",x"2B",x"D7",x"7B", -- 0x2B20
    x"C9",x"3E",x"01",x"32",x"9C",x"40",x"C1",x"CD", -- 0x2B28
    x"10",x"1B",x"C5",x"21",x"FF",x"FF",x"22",x"A2", -- 0x2B30
    x"40",x"E1",x"D1",x"4E",x"23",x"46",x"23",x"78", -- 0x2B38
    x"B1",x"CA",x"19",x"1A",x"CD",x"DF",x"41",x"CD", -- 0x2B40
    x"9B",x"1D",x"C5",x"4E",x"23",x"46",x"23",x"C5", -- 0x2B48
    x"E3",x"EB",x"DF",x"C1",x"DA",x"18",x"1A",x"E3", -- 0x2B50
    x"E5",x"C5",x"EB",x"22",x"EC",x"40",x"CD",x"AF", -- 0x2B58
    x"0F",x"3E",x"20",x"E1",x"CD",x"2A",x"03",x"CD", -- 0x2B60
    x"7E",x"2B",x"2A",x"A7",x"40",x"CD",x"75",x"2B", -- 0x2B68
    x"CD",x"FE",x"20",x"18",x"BE",x"7E",x"B7",x"C8", -- 0x2B70
    x"CD",x"2A",x"03",x"23",x"18",x"F7",x"E5",x"2A", -- 0x2B78
    x"A7",x"40",x"44",x"4D",x"E1",x"16",x"FF",x"18", -- 0x2B80
    x"03",x"03",x"15",x"C8",x"7E",x"B7",x"23",x"02", -- 0x2B88
    x"C8",x"F2",x"D2",x"3F",x"FE",x"FB",x"20",x"08", -- 0x2B90
    x"0B",x"0B",x"0B",x"0B",x"14",x"14",x"14",x"14", -- 0x2B98
    x"FE",x"95",x"CC",x"24",x"0B",x"D6",x"7F",x"E5", -- 0x2BA0
    x"5F",x"CD",x"AD",x"39",x"7E",x"B7",x"23",x"F2", -- 0x2BA8
    x"AC",x"2B",x"1D",x"20",x"F7",x"E6",x"7F",x"02", -- 0x2BB0
    x"03",x"15",x"CA",x"D8",x"28",x"7E",x"23",x"B7", -- 0x2BB8
    x"F2",x"B7",x"2B",x"E1",x"18",x"C6",x"CD",x"10", -- 0x2BC0
    x"1B",x"D1",x"C5",x"C5",x"CD",x"2C",x"1B",x"30", -- 0x2BC8
    x"05",x"54",x"5D",x"E3",x"E5",x"DF",x"D2",x"4A", -- 0x2BD0
    x"1E",x"21",x"29",x"19",x"CD",x"A7",x"28",x"C1", -- 0x2BD8
    x"21",x"E8",x"1A",x"E3",x"EB",x"2A",x"F9",x"40", -- 0x2BE0
    x"1A",x"02",x"03",x"13",x"DF",x"20",x"F9",x"60", -- 0x2BE8
    x"69",x"22",x"F9",x"40",x"C9",x"CD",x"37",x"23", -- 0x2BF0
    x"E5",x"CD",x"13",x"2A",x"F5",x"C5",x"D5",x"E5", -- 0x2BF8
    x"CD",x"3F",x"02",x"E1",x"D1",x"C1",x"F1",x"1A", -- 0x2C00
    x"CD",x"1F",x"02",x"2A",x"A4",x"40",x"EB",x"2A", -- 0x2C08
    x"F9",x"40",x"1A",x"13",x"CD",x"1F",x"02",x"DF", -- 0x2C10
    x"20",x"F8",x"00",x"00",x"00",x"E1",x"C9",x"00", -- 0x2C18
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AF", -- 0x2C20
    x"01",x"2F",x"23",x"F5",x"2B",x"D7",x"3E",x"00", -- 0x2C28
    x"28",x"07",x"CD",x"37",x"23",x"CD",x"13",x"2A", -- 0x2C30
    x"1A",x"6F",x"F1",x"B7",x"67",x"22",x"21",x"41", -- 0x2C38
    x"CC",x"4D",x"1B",x"2A",x"21",x"41",x"EB",x"F5", -- 0x2C40
    x"C5",x"D5",x"E5",x"CD",x"4C",x"02",x"E1",x"D1", -- 0x2C48
    x"C1",x"F1",x"CD",x"ED",x"01",x"1C",x"1D",x"28", -- 0x2C50
    x"03",x"BB",x"20",x"37",x"2A",x"A4",x"40",x"06", -- 0x2C58
    x"03",x"CD",x"ED",x"01",x"5F",x"96",x"A2",x"20", -- 0x2C60
    x"21",x"73",x"CD",x"6C",x"19",x"7E",x"B7",x"23", -- 0x2C68
    x"20",x"ED",x"CD",x"E4",x"01",x"10",x"EA",x"22", -- 0x2C70
    x"F9",x"40",x"21",x"29",x"19",x"CD",x"A7",x"28", -- 0x2C78
    x"00",x"00",x"00",x"2A",x"A4",x"40",x"E5",x"C3", -- 0x2C80
    x"E8",x"1A",x"21",x"A5",x"2C",x"CD",x"79",x"35", -- 0x2C88
    x"C3",x"18",x"1A",x"32",x"26",x"44",x"06",x"03", -- 0x2C90
    x"CD",x"ED",x"01",x"B7",x"20",x"F8",x"10",x"F8", -- 0x2C98
    x"00",x"00",x"00",x"18",x"A2",x"42",x"41",x"44", -- 0x2CA0
    x"0D",x"00",x"CD",x"7F",x"0A",x"7E",x"C3",x"F8", -- 0x2CA8
    x"27",x"CD",x"02",x"2B",x"D5",x"CF",x"2C",x"CD", -- 0x2CB0
    x"1C",x"2B",x"D1",x"12",x"C9",x"CD",x"38",x"23", -- 0x2CB8
    x"CD",x"F4",x"0A",x"CF",x"3B",x"EB",x"2A",x"21", -- 0x2CC0
    x"41",x"18",x"08",x"3A",x"DE",x"40",x"B7",x"28", -- 0x2CC8
    x"0C",x"D1",x"EB",x"E5",x"AF",x"32",x"DE",x"40", -- 0x2CD0
    x"BA",x"F5",x"D5",x"46",x"B0",x"CA",x"4A",x"1E", -- 0x2CD8
    x"23",x"4E",x"23",x"66",x"69",x"18",x"1C",x"58", -- 0x2CE0
    x"E5",x"0E",x"02",x"7E",x"23",x"FE",x"25",x"CA", -- 0x2CE8
    x"17",x"2E",x"FE",x"20",x"20",x"03",x"0C",x"10", -- 0x2CF0
    x"F2",x"E1",x"43",x"3E",x"25",x"CD",x"49",x"2E", -- 0x2CF8
    x"CD",x"2A",x"03",x"AF",x"5F",x"57",x"CD",x"49", -- 0x2D00
    x"2E",x"57",x"7E",x"23",x"FE",x"21",x"CA",x"14", -- 0x2D08
    x"2E",x"FE",x"23",x"28",x"37",x"05",x"CA",x"FE", -- 0x2D10
    x"2D",x"FE",x"2B",x"3E",x"08",x"28",x"E7",x"2B", -- 0x2D18
    x"7E",x"23",x"FE",x"2E",x"28",x"40",x"FE",x"25", -- 0x2D20
    x"28",x"BD",x"BE",x"20",x"D0",x"FE",x"24",x"28", -- 0x2D28
    x"14",x"FE",x"2A",x"20",x"C8",x"78",x"FE",x"02", -- 0x2D30
    x"23",x"38",x"03",x"7E",x"FE",x"24",x"3E",x"20", -- 0x2D38
    x"20",x"07",x"05",x"1C",x"FE",x"AF",x"C6",x"10", -- 0x2D40
    x"23",x"1C",x"82",x"57",x"1C",x"0E",x"00",x"05", -- 0x2D48
    x"28",x"47",x"7E",x"23",x"FE",x"2E",x"28",x"18", -- 0x2D50
    x"FE",x"23",x"28",x"F0",x"FE",x"2C",x"20",x"1A", -- 0x2D58
    x"7A",x"F6",x"40",x"57",x"18",x"E6",x"7E",x"FE", -- 0x2D60
    x"23",x"3E",x"2E",x"20",x"90",x"0E",x"01",x"23", -- 0x2D68
    x"0C",x"05",x"28",x"25",x"7E",x"23",x"FE",x"23", -- 0x2D70
    x"28",x"F6",x"D5",x"11",x"97",x"2D",x"D5",x"54", -- 0x2D78
    x"5D",x"FE",x"5B",x"C0",x"BE",x"C0",x"23",x"BE", -- 0x2D80
    x"C0",x"23",x"BE",x"C0",x"23",x"78",x"D6",x"04", -- 0x2D88
    x"D8",x"D1",x"D1",x"47",x"14",x"23",x"CA",x"EB", -- 0x2D90
    x"D1",x"7A",x"2B",x"1C",x"E6",x"08",x"20",x"15", -- 0x2D98
    x"1D",x"78",x"B7",x"28",x"10",x"7E",x"D6",x"2D", -- 0x2DA0
    x"28",x"06",x"FE",x"FE",x"20",x"07",x"3E",x"08", -- 0x2DA8
    x"C6",x"04",x"82",x"57",x"05",x"E1",x"F1",x"28", -- 0x2DB0
    x"50",x"C5",x"D5",x"CD",x"37",x"23",x"D1",x"C1", -- 0x2DB8
    x"C5",x"E5",x"43",x"78",x"81",x"FE",x"19",x"D2", -- 0x2DC0
    x"4A",x"1E",x"7A",x"F6",x"80",x"CD",x"BE",x"0F", -- 0x2DC8
    x"CD",x"A7",x"28",x"E1",x"2B",x"D7",x"37",x"28", -- 0x2DD0
    x"0D",x"32",x"DE",x"40",x"FE",x"3B",x"28",x"05", -- 0x2DD8
    x"FE",x"2C",x"C2",x"97",x"19",x"D7",x"C1",x"EB", -- 0x2DE0
    x"E1",x"E5",x"F5",x"D5",x"7E",x"90",x"23",x"4E", -- 0x2DE8
    x"23",x"66",x"69",x"16",x"00",x"5F",x"19",x"78", -- 0x2DF0
    x"B7",x"C2",x"03",x"2D",x"18",x"06",x"CD",x"49", -- 0x2DF8
    x"2E",x"CD",x"2A",x"03",x"E1",x"F1",x"C2",x"CB", -- 0x2E00
    x"2C",x"DC",x"FE",x"20",x"E3",x"CD",x"DD",x"29", -- 0x2E08
    x"E1",x"C3",x"69",x"21",x"0E",x"01",x"3E",x"F1", -- 0x2E10
    x"05",x"CD",x"49",x"2E",x"E1",x"F1",x"28",x"E9", -- 0x2E18
    x"C5",x"CD",x"37",x"23",x"CD",x"F4",x"0A",x"C1", -- 0x2E20
    x"C5",x"E5",x"2A",x"21",x"41",x"41",x"0E",x"00", -- 0x2E28
    x"C5",x"CD",x"68",x"2A",x"CD",x"AA",x"28",x"2A", -- 0x2E30
    x"21",x"41",x"F1",x"96",x"47",x"3E",x"20",x"04", -- 0x2E38
    x"05",x"CA",x"D3",x"2D",x"CD",x"2A",x"03",x"18", -- 0x2E40
    x"F7",x"F5",x"7A",x"B7",x"3E",x"2B",x"C4",x"2A", -- 0x2E48
    x"03",x"F1",x"C9",x"32",x"9A",x"40",x"2A",x"EA", -- 0x2E50
    x"40",x"B4",x"A5",x"3C",x"EB",x"C8",x"18",x"04", -- 0x2E58
    x"CD",x"4F",x"1E",x"C0",x"E1",x"EB",x"22",x"EC", -- 0x2E60
    x"40",x"EB",x"CD",x"2C",x"1B",x"D2",x"D9",x"1E", -- 0x2E68
    x"60",x"69",x"23",x"23",x"4E",x"23",x"46",x"23", -- 0x2E70
    x"C5",x"CD",x"7E",x"2B",x"E1",x"E5",x"CD",x"AF", -- 0x2E78
    x"0F",x"3E",x"20",x"CD",x"2A",x"03",x"2A",x"A7", -- 0x2E80
    x"40",x"3E",x"0E",x"CD",x"2A",x"03",x"E5",x"0E", -- 0x2E88
    x"FF",x"0C",x"7E",x"B7",x"23",x"20",x"FA",x"E1", -- 0x2E90
    x"47",x"16",x"00",x"CD",x"84",x"03",x"D6",x"30", -- 0x2E98
    x"38",x"0E",x"FE",x"0A",x"30",x"0A",x"5F",x"7A", -- 0x2EA0
    x"07",x"07",x"82",x"07",x"83",x"57",x"18",x"EB", -- 0x2EA8
    x"E5",x"21",x"99",x"2E",x"E3",x"15",x"14",x"C2", -- 0x2EB0
    x"BB",x"2E",x"14",x"FE",x"D8",x"CA",x"D2",x"2F", -- 0x2EB8
    x"FE",x"DD",x"CA",x"E0",x"2F",x"FE",x"F0",x"28", -- 0x2EC0
    x"41",x"FE",x"31",x"38",x"02",x"D6",x"20",x"FE", -- 0x2EC8
    x"21",x"CA",x"F6",x"2F",x"FE",x"1C",x"CA",x"40", -- 0x2ED0
    x"2F",x"FE",x"23",x"28",x"3F",x"FE",x"19",x"CA", -- 0x2ED8
    x"7D",x"2F",x"FE",x"14",x"CA",x"4A",x"2F",x"FE", -- 0x2EE0
    x"13",x"CA",x"65",x"2F",x"FE",x"15",x"CA",x"E3", -- 0x2EE8
    x"2F",x"FE",x"28",x"CA",x"78",x"2F",x"FE",x"1B", -- 0x2EF0
    x"28",x"1C",x"FE",x"18",x"CA",x"75",x"2F",x"FE", -- 0x2EF8
    x"11",x"C0",x"C1",x"D1",x"CD",x"FE",x"20",x"C3", -- 0x2F00
    x"65",x"2E",x"7E",x"B7",x"C8",x"04",x"CD",x"2A", -- 0x2F08
    x"03",x"23",x"15",x"20",x"F5",x"C9",x"E5",x"21", -- 0x2F10
    x"5F",x"2F",x"E3",x"37",x"F5",x"CD",x"84",x"03", -- 0x2F18
    x"5F",x"F1",x"F5",x"DC",x"5F",x"2F",x"7E",x"B7", -- 0x2F20
    x"CA",x"3E",x"2F",x"CD",x"2A",x"03",x"F1",x"F5", -- 0x2F28
    x"DC",x"A1",x"2F",x"38",x"02",x"23",x"04",x"7E", -- 0x2F30
    x"BB",x"20",x"EB",x"15",x"20",x"E8",x"F1",x"C9", -- 0x2F38
    x"CD",x"75",x"2B",x"CD",x"FE",x"20",x"C1",x"C3", -- 0x2F40
    x"7C",x"2E",x"7E",x"B7",x"C8",x"3E",x"21",x"CD", -- 0x2F48
    x"2A",x"03",x"7E",x"B7",x"28",x"09",x"CD",x"2A", -- 0x2F50
    x"03",x"CD",x"A1",x"2F",x"15",x"20",x"F3",x"3E", -- 0x2F58
    x"21",x"CD",x"2A",x"03",x"C9",x"7E",x"B7",x"C8", -- 0x2F60
    x"CD",x"84",x"03",x"77",x"CD",x"2A",x"03",x"23", -- 0x2F68
    x"04",x"15",x"20",x"F1",x"C9",x"36",x"00",x"48", -- 0x2F70
    x"16",x"FF",x"CD",x"0A",x"2F",x"CD",x"84",x"03", -- 0x2F78
    x"B7",x"CA",x"7D",x"2F",x"FE",x"08",x"28",x"0A", -- 0x2F80
    x"FE",x"0D",x"CA",x"E0",x"2F",x"FE",x"1B",x"C8", -- 0x2F88
    x"20",x"1E",x"3E",x"08",x"05",x"04",x"28",x"1F", -- 0x2F90
    x"CD",x"2A",x"03",x"2B",x"05",x"11",x"7D",x"2F", -- 0x2F98
    x"D5",x"E5",x"0D",x"7E",x"B7",x"37",x"CA",x"90", -- 0x2FA0
    x"08",x"23",x"7E",x"2B",x"77",x"23",x"18",x"F3", -- 0x2FA8
    x"F5",x"79",x"FE",x"FF",x"38",x"03",x"F1",x"18", -- 0x2FB0
    x"C4",x"90",x"0C",x"04",x"C5",x"EB",x"6F",x"26", -- 0x2FB8
    x"00",x"19",x"44",x"4D",x"23",x"CD",x"58",x"19", -- 0x2FC0
    x"C1",x"F1",x"77",x"CD",x"2A",x"03",x"23",x"C3", -- 0x2FC8
    x"7D",x"2F",x"78",x"B7",x"C8",x"05",x"2B",x"3E", -- 0x2FD0
    x"08",x"CD",x"2A",x"03",x"15",x"20",x"F3",x"C9", -- 0x2FD8
    x"CD",x"75",x"2B",x"CD",x"FE",x"20",x"C1",x"D1", -- 0x2FE0
    x"7A",x"A3",x"3C",x"2A",x"A7",x"40",x"2B",x"C8", -- 0x2FE8
    x"37",x"23",x"F5",x"C3",x"98",x"1A",x"C1",x"D1", -- 0x2FF0
    x"C3",x"19",x"1A",x"DE",x"C3",x"C3",x"44",x"B2", -- 0x2FF8
    x"C3",x"15",x"34",x"E5",x"21",x"18",x"40",x"CB", -- 0x3000
    x"7E",x"28",x"12",x"CB",x"BE",x"FE",x"31",x"38", -- 0x3008
    x"0C",x"FE",x"39",x"30",x"08",x"D6",x"31",x"CD", -- 0x3010
    x"21",x"36",x"E1",x"18",x"E3",x"E1",x"C3",x"E3", -- 0x3018
    x"05",x"FF",x"FE",x"C0",x"C3",x"05",x"31",x"D6", -- 0x3020
    x"C0",x"CA",x"08",x"31",x"47",x"3E",x"20",x"C5", -- 0x3028
    x"CD",x"84",x"31",x"C1",x"10",x"F7",x"C3",x"08", -- 0x3030
    x"31",x"23",x"E5",x"CD",x"65",x"31",x"EB",x"E1", -- 0x3038
    x"DF",x"C0",x"11",x"D8",x"FF",x"19",x"C9",x"C5", -- 0x3040
    x"E5",x"06",x"02",x"0E",x"FA",x"ED",x"79",x"0C", -- 0x3048
    x"ED",x"61",x"3C",x"65",x"10",x"F5",x"E1",x"C1", -- 0x3050
    x"C9",x"E5",x"21",x"07",x"20",x"18",x"04",x"E5", -- 0x3058
    x"2A",x"19",x"40",x"3E",x"0A",x"CD",x"47",x"30", -- 0x3060
    x"7C",x"E1",x"E5",x"D5",x"FE",x"20",x"C4",x"14", -- 0x3068
    x"36",x"00",x"3E",x"0E",x"CD",x"47",x"30",x"D1", -- 0x3070
    x"E1",x"C9",x"E5",x"D5",x"F5",x"C3",x"F8",x"35", -- 0x3078
    x"19",x"E5",x"21",x"90",x"43",x"11",x"00",x"00", -- 0x3080
    x"3A",x"23",x"40",x"5F",x"19",x"7E",x"E1",x"77", -- 0x3088
    x"F1",x"D1",x"E1",x"C9",x"03",x"01",x"02",x"04", -- 0x3090
    x"06",x"08",x"09",x"0A",x"05",x"E5",x"D5",x"C5", -- 0x3098
    x"2A",x"20",x"40",x"E5",x"CD",x"65",x"31",x"EB", -- 0x30A0
    x"E1",x"B7",x"ED",x"52",x"7D",x"C1",x"D1",x"E1", -- 0x30A8
    x"C9",x"7B",x"5F",x"3A",x"9C",x"40",x"B7",x"FA", -- 0x30B0
    x"4A",x"1E",x"28",x"05",x"3A",x"9E",x"40",x"18", -- 0x30B8
    x"03",x"3A",x"9D",x"40",x"BB",x"30",x"0B",x"C5", -- 0x30C0
    x"43",x"5F",x"78",x"C1",x"93",x"30",x"FD",x"83", -- 0x30C8
    x"5F",x"C9",x"7B",x"C9",x"21",x"E7",x"03",x"DF", -- 0x30D0
    x"E1",x"DA",x"4A",x"1E",x"C3",x"7E",x"20",x"CD", -- 0x30D8
    x"9D",x"30",x"5F",x"C9",x"DD",x"6E",x"03",x"DD", -- 0x30E0
    x"66",x"04",x"DA",x"7D",x"31",x"DD",x"7E",x"05", -- 0x30E8
    x"B7",x"20",x"05",x"CD",x"59",x"30",x"18",x"03", -- 0x30F0
    x"CD",x"5F",x"30",x"79",x"FE",x"20",x"38",x"22", -- 0x30F8
    x"FE",x"80",x"D2",x"22",x"30",x"CD",x"84",x"31", -- 0x3100
    x"7E",x"57",x"DD",x"7E",x"05",x"B7",x"28",x"08", -- 0x3108
    x"DD",x"72",x"05",x"CD",x"5F",x"30",x"18",x"03", -- 0x3110
    x"CD",x"59",x"30",x"DD",x"75",x"03",x"DD",x"74", -- 0x3118
    x"04",x"C9",x"11",x"08",x"31",x"D5",x"FE",x"08", -- 0x3120
    x"CA",x"DF",x"31",x"FE",x"0A",x"D8",x"FE",x"0E", -- 0x3128
    x"DA",x"C9",x"31",x"CA",x"F8",x"31",x"FE",x"0F", -- 0x3130
    x"CA",x"FD",x"31",x"FE",x"18",x"D8",x"FE",x"18", -- 0x3138
    x"CA",x"E5",x"31",x"FE",x"19",x"CA",x"39",x"30", -- 0x3140
    x"FE",x"1A",x"CA",x"00",x"32",x"FE",x"1B",x"CA", -- 0x3148
    x"12",x"32",x"FE",x"1C",x"CA",x"D4",x"31",x"FE", -- 0x3150
    x"1D",x"CA",x"D9",x"31",x"FE",x"1E",x"28",x"5F", -- 0x3158
    x"FE",x"1F",x"28",x"45",x"C9",x"11",x"00",x"BC", -- 0x3160
    x"06",x"01",x"19",x"11",x"28",x"00",x"B7",x"ED", -- 0x3168
    x"52",x"38",x"03",x"04",x"18",x"F5",x"21",x"D8", -- 0x3170
    x"43",x"19",x"10",x"FD",x"C9",x"DD",x"7E",x"05", -- 0x3178
    x"B7",x"C0",x"7E",x"C9",x"CD",x"7A",x"30",x"77", -- 0x3180
    x"23",x"11",x"E8",x"47",x"DF",x"D8",x"21",x"E8", -- 0x3188
    x"47",x"11",x"D8",x"FF",x"19",x"E5",x"CD",x"39", -- 0x3190
    x"36",x"ED",x"A0",x"D9",x"ED",x"A0",x"D9",x"78", -- 0x3198
    x"B1",x"20",x"F6",x"D9",x"E1",x"D1",x"C1",x"D9", -- 0x31A0
    x"E1",x"11",x"E8",x"47",x"E5",x"CD",x"E0",x"31", -- 0x31A8
    x"23",x"DF",x"20",x"F9",x"E1",x"C9",x"FD",x"E5", -- 0x31B0
    x"18",x"68",x"FD",x"E1",x"C3",x"83",x"2C",x"E5", -- 0x31B8
    x"CD",x"65",x"31",x"EB",x"19",x"EB",x"E1",x"18", -- 0x31C0
    x"E3",x"CD",x"1B",x"36",x"19",x"11",x"E8",x"47", -- 0x31C8
    x"DF",x"28",x"BE",x"C9",x"21",x"00",x"44",x"18", -- 0x31D0
    x"03",x"CD",x"65",x"31",x"C3",x"5F",x"30",x"2B", -- 0x31D8
    x"3E",x"20",x"C3",x"EE",x"35",x"E5",x"CD",x"65", -- 0x31E0
    x"31",x"EB",x"E1",x"DF",x"28",x"03",x"2B",x"18", -- 0x31E8
    x"EB",x"2B",x"11",x"28",x"00",x"19",x"18",x"E4", -- 0x31F0
    x"7E",x"DD",x"77",x"05",x"C9",x"AF",x"18",x"F9", -- 0x31F8
    x"CD",x"07",x"36",x"19",x"B7",x"3F",x"11",x"E8", -- 0x3200
    x"47",x"DF",x"38",x"04",x"11",x"40",x"FC",x"19", -- 0x3208
    x"18",x"CA",x"CD",x"0F",x"36",x"19",x"11",x"00", -- 0x3210
    x"44",x"DF",x"30",x"04",x"11",x"E8",x"03",x"19", -- 0x3218
    x"18",x"BA",x"2B",x"D7",x"20",x"06",x"11",x"0A", -- 0x3220
    x"00",x"D5",x"18",x"13",x"D2",x"4A",x"1E",x"CD", -- 0x3228
    x"5A",x"1E",x"CF",x"2C",x"30",x"F6",x"D5",x"CD", -- 0x3230
    x"5A",x"1E",x"7A",x"B3",x"CA",x"4A",x"1E",x"ED", -- 0x3238
    x"53",x"E4",x"40",x"D1",x"ED",x"53",x"E2",x"40", -- 0x3240
    x"FD",x"2A",x"F9",x"40",x"11",x"00",x"01",x"FD", -- 0x3248
    x"19",x"FD",x"E5",x"2A",x"A4",x"40",x"E5",x"7E", -- 0x3250
    x"23",x"B6",x"28",x"4A",x"23",x"23",x"CD",x"BA", -- 0x3258
    x"33",x"23",x"28",x"F3",x"CD",x"D8",x"33",x"2B", -- 0x3260
    x"28",x"F4",x"23",x"E5",x"D5",x"FD",x"E5",x"D1", -- 0x3268
    x"2A",x"B1",x"40",x"ED",x"52",x"DA",x"7A",x"19", -- 0x3270
    x"11",x"04",x"00",x"ED",x"52",x"DA",x"7A",x"19", -- 0x3278
    x"FD",x"70",x"00",x"E1",x"CD",x"5A",x"1E",x"FD", -- 0x3280
    x"73",x"01",x"FD",x"72",x"02",x"FD",x"36",x"03", -- 0x3288
    x"00",x"CD",x"B1",x"33",x"E1",x"2B",x"23",x"7E", -- 0x3290
    x"FE",x"20",x"28",x"FA",x"FE",x"2C",x"28",x"03", -- 0x3298
    x"2B",x"18",x"BB",x"23",x"18",x"BE",x"FD",x"36", -- 0x32A0
    x"00",x"FF",x"E1",x"FD",x"E1",x"ED",x"5B",x"E2", -- 0x32A8
    x"40",x"D5",x"FD",x"E5",x"E5",x"D5",x"CD",x"C2", -- 0x32B0
    x"09",x"7A",x"B3",x"28",x"41",x"EB",x"D1",x"FD", -- 0x32B8
    x"E5",x"FD",x"7E",x"00",x"3C",x"28",x"21",x"FD", -- 0x32C0
    x"7E",x"03",x"B7",x"20",x"16",x"FD",x"7E",x"01", -- 0x32C8
    x"B9",x"20",x"10",x"FD",x"7E",x"02",x"B8",x"20", -- 0x32D0
    x"0A",x"FD",x"73",x"01",x"FD",x"72",x"02",x"FD", -- 0x32D8
    x"36",x"03",x"01",x"CD",x"B1",x"33",x"18",x"D9", -- 0x32E0
    x"FD",x"E1",x"E5",x"2A",x"E4",x"40",x"19",x"DA", -- 0x32E8
    x"7A",x"19",x"EB",x"21",x"F8",x"FF",x"ED",x"52", -- 0x32F0
    x"DA",x"7A",x"19",x"E1",x"18",x"B7",x"D1",x"E1", -- 0x32F8
    x"FD",x"E1",x"D1",x"7E",x"23",x"B6",x"CA",x"BA", -- 0x3300
    x"31",x"23",x"73",x"23",x"72",x"CD",x"BA",x"33", -- 0x3308
    x"23",x"20",x"09",x"E5",x"2A",x"E4",x"40",x"19", -- 0x3310
    x"EB",x"E1",x"18",x"E7",x"E5",x"D5",x"CD",x"D8", -- 0x3318
    x"33",x"D1",x"E1",x"2B",x"28",x"E7",x"23",x"7E", -- 0x3320
    x"FE",x"20",x"28",x"FA",x"D5",x"E5",x"FD",x"6E", -- 0x3328
    x"01",x"FD",x"66",x"02",x"CD",x"94",x"33",x"FD", -- 0x3330
    x"4E",x"00",x"CD",x"B1",x"33",x"EB",x"E1",x"CD", -- 0x3338
    x"F8",x"33",x"D1",x"2B",x"23",x"7E",x"FE",x"20", -- 0x3340
    x"28",x"FA",x"FE",x"2C",x"28",x"03",x"2B",x"18", -- 0x3348
    x"BC",x"23",x"18",x"C8",x"D5",x"C5",x"E5",x"E5", -- 0x3350
    x"D1",x"D5",x"D5",x"2A",x"F9",x"40",x"E5",x"2B", -- 0x3358
    x"13",x"10",x"FC",x"22",x"F9",x"40",x"E1",x"C1", -- 0x3360
    x"ED",x"42",x"23",x"E5",x"C1",x"E1",x"EB",x"ED", -- 0x3368
    x"B0",x"E1",x"C1",x"D1",x"C9",x"D5",x"C5",x"E5", -- 0x3370
    x"2A",x"F9",x"40",x"E5",x"D1",x"23",x"10",x"FD", -- 0x3378
    x"22",x"F9",x"40",x"C1",x"C5",x"E5",x"B7",x"ED", -- 0x3380
    x"42",x"E5",x"C1",x"03",x"E1",x"EB",x"ED",x"B8", -- 0x3388
    x"E1",x"C1",x"D1",x"C9",x"D5",x"22",x"21",x"41", -- 0x3390
    x"01",x"00",x"00",x"2A",x"A7",x"40",x"E5",x"CD", -- 0x3398
    x"2F",x"13",x"E1",x"06",x"05",x"7E",x"D6",x"30", -- 0x33A0
    x"20",x"05",x"23",x"10",x"F8",x"2B",x"04",x"D1", -- 0x33A8
    x"C9",x"FD",x"23",x"FD",x"23",x"FD",x"23",x"FD", -- 0x33B0
    x"23",x"C9",x"23",x"7E",x"B7",x"C8",x"FE",x"8D", -- 0x33B8
    x"28",x"0C",x"FE",x"91",x"28",x"08",x"FE",x"CA", -- 0x33C0
    x"28",x"04",x"FE",x"95",x"20",x"EC",x"2B",x"7E", -- 0x33C8
    x"FE",x"FF",x"23",x"7E",x"28",x"E4",x"A7",x"C9", -- 0x33D0
    x"ED",x"5B",x"A7",x"40",x"D5",x"06",x"00",x"7E", -- 0x33D8
    x"FE",x"20",x"28",x"0B",x"FE",x"30",x"38",x"0A", -- 0x33E0
    x"FE",x"3A",x"30",x"06",x"04",x"12",x"13",x"23", -- 0x33E8
    x"18",x"ED",x"AF",x"12",x"D1",x"04",x"05",x"C9", -- 0x33F0
    x"C5",x"78",x"99",x"28",x"10",x"05",x"28",x"08", -- 0x33F8
    x"0D",x"20",x"F6",x"CD",x"75",x"33",x"18",x"05", -- 0x3400
    x"41",x"05",x"CD",x"54",x"33",x"C1",x"1A",x"77", -- 0x3408
    x"13",x"23",x"10",x"FA",x"C9",x"CD",x"49",x"00", -- 0x3410
    x"FE",x"5C",x"38",x"3C",x"FE",x"60",x"30",x"38", -- 0x3418
    x"D6",x"5B",x"57",x"78",x"FE",x"07",x"38",x"ED", -- 0x3420
    x"7A",x"C5",x"E5",x"21",x"49",x"43",x"11",x"07", -- 0x3428
    x"00",x"19",x"3D",x"20",x"FC",x"D1",x"06",x"07", -- 0x3430
    x"7E",x"FE",x"00",x"28",x"12",x"12",x"D5",x"CD", -- 0x3438
    x"33",x"00",x"D1",x"23",x"13",x"10",x"F1",x"EB", -- 0x3440
    x"C1",x"78",x"D6",x"07",x"47",x"18",x"C6",x"EB", -- 0x3448
    x"78",x"C1",x"80",x"D6",x"07",x"47",x"3E",x"0D", -- 0x3450
    x"FE",x"7C",x"DA",x"03",x"30",x"FE",x"80",x"D2", -- 0x3458
    x"03",x"30",x"D6",x"77",x"18",x"BC",x"2B",x"D7", -- 0x3460
    x"D2",x"4A",x"1E",x"D6",x"30",x"F5",x"23",x"CF", -- 0x3468
    x"D5",x"CF",x"22",x"F1",x"FE",x"01",x"DA",x"4A", -- 0x3470
    x"1E",x"FE",x"09",x"30",x"EB",x"E5",x"21",x"49", -- 0x3478
    x"43",x"11",x"07",x"00",x"19",x"3D",x"20",x"FC", -- 0x3480
    x"EB",x"E1",x"2B",x"06",x"07",x"D7",x"FE",x"22", -- 0x3488
    x"28",x"0C",x"FE",x"00",x"28",x"0A",x"12",x"13", -- 0x3490
    x"10",x"F3",x"23",x"CF",x"22",x"C9",x"3E",x"20", -- 0x3498
    x"12",x"05",x"28",x"03",x"13",x"18",x"F9",x"B7", -- 0x34A0
    x"C8",x"18",x"F0",x"4C",x"49",x"53",x"54",x"20", -- 0x34A8
    x"20",x"20",x"52",x"55",x"4E",x"20",x"20",x"20", -- 0x34B0
    x"20",x"41",x"55",x"54",x"4F",x"20",x"20",x"20", -- 0x34B8
    x"45",x"44",x"49",x"54",x"20",x"20",x"20",x"52", -- 0x34C0
    x"45",x"4E",x"55",x"4D",x"20",x"20",x"53",x"59", -- 0x34C8
    x"53",x"54",x"45",x"4D",x"00",x"43",x"4C",x"4F", -- 0x34D0
    x"41",x"44",x"20",x"20",x"43",x"53",x"41",x"56", -- 0x34D8
    x"45",x"20",x"22",x"D7",x"FE",x"48",x"11",x"00", -- 0x34E0
    x"00",x"20",x"3D",x"23",x"CD",x"16",x"35",x"DA", -- 0x34E8
    x"97",x"19",x"CD",x"FE",x"34",x"E5",x"EB",x"CD", -- 0x34F0
    x"9A",x"0A",x"E1",x"2B",x"D7",x"C9",x"CD",x"16", -- 0x34F8
    x"35",x"D8",x"06",x"04",x"CD",x"09",x"35",x"18", -- 0x3500
    x"F5",x"CB",x"23",x"CB",x"12",x"DA",x"B2",x"07", -- 0x3508
    x"10",x"F7",x"B3",x"5F",x"23",x"C9",x"CD",x"3D", -- 0x3510
    x"1E",x"38",x"06",x"D6",x"37",x"FE",x"10",x"3F", -- 0x3518
    x"C9",x"D6",x"30",x"D8",x"FE",x"0A",x"3F",x"C9", -- 0x3520
    x"FE",x"4F",x"C2",x"97",x"19",x"23",x"CD",x"41", -- 0x3528
    x"35",x"DA",x"97",x"19",x"CD",x"41",x"35",x"DA", -- 0x3530
    x"F5",x"34",x"06",x"03",x"CD",x"09",x"35",x"18", -- 0x3538
    x"F3",x"7E",x"D6",x"30",x"D8",x"FE",x"08",x"3F", -- 0x3540
    x"C9",x"2B",x"AF",x"1E",x"D9",x"C3",x"29",x"2C", -- 0x3548
    x"11",x"00",x"00",x"CD",x"16",x"35",x"DA",x"97", -- 0x3550
    x"19",x"C9",x"CD",x"50",x"35",x"CD",x"FE",x"34", -- 0x3558
    x"E5",x"EB",x"11",x"67",x"35",x"D5",x"E9",x"E1", -- 0x3560
    x"C9",x"03",x"05",x"02",x"04",x"06",x"08",x"01", -- 0x3568
    x"0E",x"09",x"10",x"07",x"0B",x"0C",x"0D",x"0A", -- 0x3570
    x"0F",x"CD",x"A7",x"28",x"11",x"09",x"00",x"D5", -- 0x3578
    x"11",x"00",x"08",x"D5",x"11",x"3E",x"10",x"D5", -- 0x3580
    x"11",x"78",x"00",x"3E",x"01",x"CD",x"2A",x"3E", -- 0x3588
    x"D1",x"3E",x"08",x"CD",x"2A",x"3E",x"D1",x"3E", -- 0x3590
    x"0C",x"CD",x"2A",x"3E",x"D1",x"3E",x"0D",x"C3", -- 0x3598
    x"32",x"3E",x"2A",x"B1",x"40",x"23",x"C3",x"F5", -- 0x35A0
    x"3C",x"CD",x"B5",x"35",x"C3",x"3F",x"02",x"CD", -- 0x35A8
    x"B5",x"35",x"C3",x"4C",x"02",x"AF",x"CD",x"01", -- 0x35B0
    x"2B",x"CF",x"2C",x"7B",x"A2",x"C6",x"02",x"D2", -- 0x35B8
    x"4A",x"1E",x"C9",x"2B",x"D7",x"28",x"1A",x"CD", -- 0x35C0
    x"1C",x"2B",x"06",x"08",x"FE",x"01",x"28",x"0B", -- 0x35C8
    x"04",x"FE",x"02",x"28",x"06",x"04",x"FE",x"03", -- 0x35D0
    x"C2",x"4A",x"1E",x"78",x"1E",x"00",x"C3",x"32", -- 0x35D8
    x"3E",x"3E",x"0A",x"11",x"00",x"00",x"CD",x"2A", -- 0x35E0
    x"3E",x"3E",x"08",x"C3",x"32",x"3E",x"77",x"CD", -- 0x35E8
    x"7A",x"30",x"23",x"CD",x"7A",x"30",x"2B",x"C9", -- 0x35F0
    x"11",x"00",x"AC",x"FE",x"20",x"C2",x"80",x"30", -- 0x35F8
    x"3A",x"90",x"43",x"19",x"C3",x"8F",x"30",x"11", -- 0x3600
    x"28",x"00",x"3E",x"20",x"C3",x"7A",x"30",x"11", -- 0x3608
    x"D8",x"FF",x"18",x"F6",x"20",x"02",x"3E",x"20", -- 0x3610
    x"C3",x"7A",x"30",x"CD",x"0A",x"36",x"C3",x"65", -- 0x3618
    x"31",x"32",x"23",x"40",x"2A",x"20",x"40",x"C3", -- 0x3620
    x"5F",x"30",x"E5",x"EB",x"11",x"28",x"00",x"19", -- 0x3628
    x"B7",x"ED",x"52",x"30",x"FC",x"19",x"7D",x"E1", -- 0x3630
    x"C9",x"D9",x"F1",x"C5",x"D5",x"E5",x"11",x"00", -- 0x3638
    x"F0",x"21",x"28",x"F0",x"01",x"C0",x"03",x"C5", -- 0x3640
    x"D9",x"11",x"00",x"44",x"21",x"28",x"44",x"C1", -- 0x3648
    x"F5",x"C9",x"7E",x"23",x"FE",x"DB",x"CA",x"C5", -- 0x3650
    x"36",x"FE",x"A0",x"CA",x"B3",x"36",x"C3",x"97", -- 0x3658
    x"19",x"3A",x"23",x"40",x"3C",x"CA",x"0D",x"37", -- 0x3660
    x"B8",x"77",x"2A",x"A4",x"40",x"2B",x"06",x"03", -- 0x3668
    x"E5",x"26",x"0F",x"CD",x"BB",x"3A",x"CB",x"57", -- 0x3670
    x"28",x"F9",x"CD",x"BB",x"3A",x"CB",x"57",x"20", -- 0x3678
    x"F9",x"26",x"0E",x"CD",x"BB",x"3A",x"E1",x"77", -- 0x3680
    x"B7",x"23",x"20",x"E2",x"10",x"E2",x"C9",x"2A", -- 0x3688
    x"A4",x"40",x"2B",x"ED",x"5B",x"F9",x"40",x"7E", -- 0x3690
    x"E5",x"6F",x"26",x"0E",x"CD",x"B2",x"3A",x"24", -- 0x3698
    x"3E",x"04",x"CD",x"B2",x"3A",x"06",x"0A",x"10", -- 0x36A0
    x"FE",x"AF",x"CD",x"B2",x"3A",x"E1",x"23",x"DF", -- 0x36A8
    x"20",x"E5",x"C9",x"E5",x"26",x"07",x"CD",x"BB", -- 0x36B0
    x"3A",x"E6",x"3F",x"F6",x"C0",x"CD",x"B2",x"3A", -- 0x36B8
    x"CD",x"8F",x"36",x"E1",x"C9",x"3E",x"07",x"D3", -- 0x36C0
    x"F8",x"3E",x"3F",x"D3",x"F9",x"CD",x"6A",x"36", -- 0x36C8
    x"C3",x"77",x"2C",x"CD",x"0D",x"26",x"D5",x"3A", -- 0x36D0
    x"AF",x"40",x"F5",x"CF",x"2C",x"CD",x"0D",x"26", -- 0x36D8
    x"C1",x"3A",x"AF",x"40",x"B8",x"C2",x"4A",x"1E", -- 0x36E0
    x"E3",x"4E",x"1A",x"77",x"79",x"12",x"23",x"13", -- 0x36E8
    x"10",x"F7",x"E1",x"C9",x"CF",x"28",x"CD",x"1C", -- 0x36F0
    x"2B",x"F5",x"CF",x"29",x"F1",x"FE",x"10",x"D2", -- 0x36F8
    x"4A",x"1E",x"E5",x"67",x"CD",x"BB",x"3A",x"C3", -- 0x3700
    x"72",x"3F",x"3A",x"14",x"43",x"E5",x"C3",x"72", -- 0x3708
    x"3F",x"10",x"0D",x"0E",x"04",x"06",x"03",x"01", -- 0x3710
    x"02",x"05",x"07",x"08",x"09",x"0A",x"0B",x"0C", -- 0x3718
    x"0F",x"10",x"0D",x"06",x"04",x"0F",x"03",x"09", -- 0x3720
    x"02",x"01",x"05",x"07",x"08",x"0A",x"0B",x"0C", -- 0x3728
    x"0E",x"10",x"05",x"02",x"04",x"0E",x"09",x"01", -- 0x3730
    x"0A",x"07",x"06",x"0D",x"03",x"08",x"0B",x"0C", -- 0x3738
    x"0F",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3740
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3748
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3750
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3758
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3760
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3768
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3770
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3778
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3780
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3788
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3790
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x3798
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37A0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37A8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37B0
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37B8
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF", -- 0x37C0
    x"FF",x"FF",x"FF",x"D5",x"11",x"1D",x"40",x"18", -- 0x37C8
    x"04",x"D5",x"11",x"25",x"40",x"E5",x"7E",x"FE", -- 0x37D0
    x"03",x"28",x"09",x"CD",x"1B",x"00",x"7E",x"FE", -- 0x37D8
    x"0D",x"23",x"20",x"F2",x"E1",x"D1",x"C9",x"7A", -- 0x37E0
    x"CD",x"EC",x"37",x"7B",x"F5",x"0F",x"0F",x"0F", -- 0x37E8
    x"0F",x"CD",x"F5",x"37",x"F1",x"E6",x"0F",x"C6", -- 0x37F0
    x"90",x"27",x"CE",x"40",x"27",x"77",x"23",x"C9", -- 0x37F8
    x"01",x"00",x"00",x"04",x"07",x"C4",x"07",x"A0", -- 0x3800
    x"1F",x"19",x"00",x"26",x"96",x"34",x"28",x"46", -- 0x3808
    x"00",x"00",x"00",x"08",x"00",x"20",x"01",x"20", -- 0x3810
    x"74",x"66",x"1F",x"7E",x"96",x"34",x"28",x"46", -- 0x3818
    x"46",x"4B",x"69",x"01",x"00",x"00",x"04",x"07", -- 0x3820
    x"C4",x"07",x"A0",x"1B",x"19",x"06",x"1F",x"34", -- 0x3828
    x"2E",x"28",x"38",x"00",x"00",x"00",x"08",x"00", -- 0x3830
    x"20",x"01",x"20",x"6E",x"66",x"08",x"7F",x"34", -- 0x3838
    x"2E",x"28",x"38",x"4C",x"51",x"71",x"3E",x"00", -- 0x3840
    x"18",x"08",x"C4",x"C2",x"3F",x"FE",x"04",x"D2", -- 0x3848
    x"4A",x"1E",x"4F",x"06",x"03",x"07",x"07",x"B1", -- 0x3850
    x"10",x"FB",x"4F",x"E5",x"2A",x"A4",x"40",x"11", -- 0x3858
    x"01",x"48",x"DF",x"28",x"09",x"21",x"00",x"48", -- 0x3860
    x"71",x"01",x"FF",x"0F",x"ED",x"B0",x"E1",x"C9", -- 0x3868
    x"3A",x"1C",x"43",x"E5",x"21",x"F0",x"42",x"CB", -- 0x3870
    x"6F",x"28",x"03",x"21",x"00",x"43",x"D3",x"FF", -- 0x3878
    x"32",x"1C",x"43",x"06",x"10",x"0E",x"FA",x"05", -- 0x3880
    x"ED",x"41",x"04",x"0C",x"ED",x"A3",x"20",x"F5", -- 0x3888
    x"E1",x"C9",x"D9",x"3A",x"1C",x"43",x"E6",x"DB", -- 0x3890
    x"CD",x"73",x"38",x"D9",x"CD",x"A7",x"28",x"C9", -- 0x3898
    x"D9",x"CD",x"70",x"38",x"D9",x"22",x"A2",x"40", -- 0x38A0
    x"C9",x"3A",x"1C",x"43",x"CB",x"EF",x"18",x"C3", -- 0x38A8
    x"3A",x"1C",x"43",x"CB",x"AF",x"18",x"BC",x"06", -- 0x38B0
    x"04",x"18",x"02",x"06",x"00",x"3A",x"1C",x"43", -- 0x38B8
    x"E6",x"FB",x"B0",x"32",x"1C",x"43",x"D3",x"FF", -- 0x38C0
    x"C9",x"CD",x"C2",x"3F",x"FE",x"10",x"D2",x"4A", -- 0x38C8
    x"1E",x"32",x"23",x"40",x"C9",x"CF",x"52",x"CD", -- 0x38D0
    x"C2",x"3F",x"FE",x"04",x"30",x"F0",x"32",x"13", -- 0x38D8
    x"43",x"C9",x"E6",x"7F",x"C0",x"EB",x"11",x"2F", -- 0x38E0
    x"39",x"C5",x"06",x"7F",x"7E",x"FE",x"61",x"38", -- 0x38E8
    x"06",x"FE",x"7B",x"30",x"02",x"E6",x"5F",x"4E", -- 0x38F0
    x"EB",x"23",x"B6",x"F2",x"F9",x"38",x"04",x"7E", -- 0x38F8
    x"E6",x"7F",x"28",x"29",x"B9",x"20",x"F2",x"EB", -- 0x3900
    x"E5",x"13",x"1A",x"B7",x"FA",x"1E",x"39",x"4F", -- 0x3908
    x"23",x"7E",x"FE",x"61",x"38",x"02",x"E6",x"5F", -- 0x3910
    x"B9",x"28",x"EE",x"E1",x"18",x"D9",x"F1",x"F1", -- 0x3918
    x"F1",x"D1",x"D1",x"E3",x"36",x"FF",x"78",x"42", -- 0x3920
    x"4B",x"D1",x"C3",x"57",x"3D",x"C1",x"F1",x"C9", -- 0x3928
    x"C3",x"4F",x"4C",x"4F",x"55",x"52",x"C6",x"43", -- 0x3930
    x"4F",x"4C",x"4F",x"55",x"CB",x"45",x"59",x"50", -- 0x3938
    x"41",x"44",x"CA",x"4F",x"59",x"D0",x"4C",x"4F", -- 0x3940
    x"54",x"C6",x"47",x"52",x"CC",x"47",x"52",x"C6", -- 0x3948
    x"43",x"4C",x"53",x"D0",x"4C",x"41",x"59",x"C3", -- 0x3950
    x"49",x"52",x"43",x"4C",x"45",x"D3",x"43",x"41", -- 0x3958
    x"4C",x"45",x"D3",x"48",x"41",x"50",x"45",x"CE", -- 0x3960
    x"53",x"48",x"41",x"50",x"45",x"D8",x"53",x"48", -- 0x3968
    x"41",x"50",x"45",x"D0",x"41",x"49",x"4E",x"54", -- 0x3970
    x"C3",x"50",x"4F",x"49",x"4E",x"54",x"CE",x"50", -- 0x3978
    x"4C",x"4F",x"54",x"D3",x"4F",x"55",x"4E",x"44", -- 0x3980
    x"C3",x"48",x"41",x"52",x"D2",x"45",x"4E",x"55", -- 0x3988
    x"4D",x"D3",x"57",x"41",x"50",x"C6",x"4B",x"45", -- 0x3990
    x"59",x"C3",x"41",x"4C",x"4C",x"D6",x"45",x"52", -- 0x3998
    x"49",x"46",x"59",x"C2",x"47",x"52",x"44",x"CE", -- 0x39A0
    x"42",x"47",x"52",x"44",x"80",x"FE",x"80",x"21", -- 0x39A8
    x"50",x"16",x"C0",x"E1",x"E3",x"7E",x"D6",x"7F", -- 0x39B0
    x"5F",x"23",x"E3",x"E5",x"2A",x"8C",x"43",x"C9", -- 0x39B8
    x"FE",x"7F",x"28",x"08",x"FE",x"3C",x"D2",x"E7", -- 0x39C0
    x"2A",x"C3",x"6A",x"1D",x"23",x"7E",x"D6",x"80", -- 0x39C8
    x"07",x"4F",x"06",x"00",x"EB",x"2A",x"8E",x"43", -- 0x39D0
    x"C3",x"72",x"1D",x"C9",x"38",x"D5",x"38",x"97", -- 0x39D8
    x"19",x"52",x"36",x"C1",x"3B",x"A9",x"38",x"B0", -- 0x39E0
    x"38",x"83",x"3C",x"61",x"3D",x"F8",x"3A",x"F1", -- 0x39E8
    x"3A",x"DD",x"3C",x"D8",x"3C",x"D3",x"3C",x"38", -- 0x39F0
    x"3E",x"97",x"19",x"BE",x"3B",x"95",x"3F",x"A8", -- 0x39F8
    x"3F",x"B6",x"31",x"D3",x"36",x"66",x"34",x"5A", -- 0x3A00
    x"35",x"49",x"35",x"E4",x"3F",x"BB",x"38",x"7E", -- 0x3A08
    x"23",x"E5",x"FE",x"31",x"CA",x"D8",x"3A",x"FE", -- 0x3A10
    x"32",x"CA",x"DC",x"3A",x"C3",x"C3",x"3A",x"7E", -- 0x3A18
    x"FE",x"28",x"28",x"26",x"16",x"04",x"FE",x"32", -- 0x3A20
    x"28",x"07",x"CB",x"3A",x"FE",x"31",x"C2",x"97", -- 0x3A28
    x"19",x"D7",x"FE",x"59",x"28",x"05",x"15",x"FE", -- 0x3A30
    x"58",x"20",x"F3",x"23",x"E5",x"CD",x"5E",x"3A", -- 0x3A38
    x"E6",x"3F",x"3C",x"18",x"16",x"18",x"F4",x"00", -- 0x3A40
    x"00",x"00",x"23",x"CD",x"1C",x"2B",x"FE",x"08", -- 0x3A48
    x"D2",x"4A",x"1E",x"57",x"CF",x"29",x"14",x"E5", -- 0x3A50
    x"CD",x"5E",x"3A",x"C3",x"72",x"3F",x"CD",x"A9", -- 0x3A58
    x"3A",x"AF",x"1E",x"80",x"B3",x"6F",x"26",x"0E", -- 0x3A60
    x"CD",x"B3",x"3A",x"24",x"CD",x"BB",x"3A",x"D5", -- 0x3A68
    x"17",x"15",x"20",x"FC",x"D1",x"7D",x"38",x"03", -- 0x3A70
    x"7B",x"2F",x"A5",x"CB",x"3B",x"30",x"E5",x"C9", -- 0x3A78
    x"C3",x"14",x"3F",x"00",x"C3",x"18",x"3F",x"CD", -- 0x3A80
    x"A9",x"3A",x"1E",x"E4",x"06",x"03",x"6A",x"26", -- 0x3A88
    x"0E",x"CD",x"B3",x"3A",x"24",x"CD",x"BB",x"3A", -- 0x3A90
    x"0E",x"04",x"1F",x"30",x"08",x"1C",x"0D",x"20", -- 0x3A98
    x"F9",x"CB",x"02",x"10",x"E9",x"16",x"3A",x"1A", -- 0x3AA0
    x"C9",x"26",x"07",x"CD",x"BB",x"3A",x"E6",x"3F", -- 0x3AA8
    x"F6",x"40",x"6F",x"0E",x"F8",x"ED",x"61",x"0C", -- 0x3AB0
    x"ED",x"69",x"C9",x"0E",x"F8",x"ED",x"61",x"0C", -- 0x3AB8
    x"ED",x"78",x"C9",x"E1",x"2B",x"CF",x"28",x"CD", -- 0x3AC0
    x"C2",x"3F",x"FE",x"02",x"D2",x"4A",x"1E",x"F5", -- 0x3AC8
    x"CF",x"29",x"F1",x"E5",x"FE",x"01",x"28",x"04", -- 0x3AD0
    x"16",x"FE",x"18",x"02",x"16",x"F7",x"CD",x"87", -- 0x3AD8
    x"3A",x"C3",x"72",x"3F",x"03",x"06",x"09",x"0C", -- 0x3AE0
    x"02",x"05",x"08",x"0A",x"01",x"04",x"07",x"0B", -- 0x3AE8
    x"00",x"CD",x"1C",x"2B",x"32",x"14",x"43",x"C9", -- 0x3AF0
    x"CD",x"1C",x"2B",x"F5",x"CF",x"2C",x"CD",x"1C", -- 0x3AF8
    x"2B",x"F5",x"CF",x"2C",x"CD",x"1C",x"2B",x"D1", -- 0x3B00
    x"C1",x"4A",x"E5",x"57",x"1E",x"00",x"26",x"80", -- 0x3B08
    x"FA",x"52",x"3B",x"CD",x"7A",x"3B",x"CD",x"7A", -- 0x3B10
    x"3B",x"CD",x"5E",x"3B",x"C5",x"D5",x"E5",x"2E", -- 0x3B18
    x"80",x"63",x"06",x"08",x"1E",x"00",x"29",x"ED", -- 0x3B20
    x"52",x"38",x"03",x"23",x"18",x"01",x"19",x"10", -- 0x3B28
    x"F5",x"7D",x"E1",x"D1",x"C1",x"84",x"67",x"7A", -- 0x3B30
    x"2E",x"00",x"9D",x"57",x"1C",x"7A",x"BB",x"C3", -- 0x3B38
    x"10",x"3B",x"C5",x"D5",x"E5",x"7B",x"80",x"6F", -- 0x3B40
    x"7A",x"81",x"67",x"CD",x"8A",x"3B",x"E1",x"D1", -- 0x3B48
    x"C1",x"C9",x"E1",x"C9",x"7B",x"ED",x"44",x"5F", -- 0x3B50
    x"C9",x"7A",x"ED",x"44",x"57",x"C9",x"CD",x"54", -- 0x3B58
    x"3B",x"CD",x"59",x"3B",x"C9",x"CD",x"54",x"3B", -- 0x3B60
    x"CD",x"42",x"3B",x"C9",x"CD",x"59",x"3B",x"CD", -- 0x3B68
    x"42",x"3B",x"C9",x"7B",x"6F",x"7A",x"5F",x"7D", -- 0x3B70
    x"57",x"C9",x"CD",x"42",x"3B",x"CD",x"65",x"3B", -- 0x3B78
    x"CD",x"6C",x"3B",x"CD",x"65",x"3B",x"CD",x"73", -- 0x3B80
    x"3B",x"C9",x"3A",x"13",x"43",x"E6",x"03",x"4F", -- 0x3B88
    x"3E",x"9F",x"BD",x"D8",x"3E",x"65",x"BC",x"D8", -- 0x3B90
    x"7D",x"6C",x"26",x"00",x"54",x"5D",x"29",x"29", -- 0x3B98
    x"19",x"29",x"29",x"29",x"5F",x"CB",x"3B",x"CB", -- 0x3BA0
    x"3B",x"16",x"48",x"19",x"E6",x"03",x"3C",x"47", -- 0x3BA8
    x"3E",x"FC",x"0F",x"0F",x"CB",x"09",x"CB",x"09", -- 0x3BB0
    x"10",x"F8",x"A6",x"B1",x"77",x"C9",x"06",x"00", -- 0x3BB8
    x"3A",x"06",x"03",x"3A",x"13",x"43",x"F5",x"A0", -- 0x3BC0
    x"32",x"13",x"43",x"CD",x"7B",x"3C",x"38",x"2F", -- 0x3BC8
    x"3A",x"15",x"43",x"F5",x"3A",x"16",x"43",x"F5", -- 0x3BD0
    x"CD",x"1C",x"2B",x"32",x"15",x"43",x"F5",x"CF", -- 0x3BD8
    x"2C",x"CD",x"1C",x"2B",x"32",x"16",x"43",x"D9", -- 0x3BE0
    x"6F",x"D1",x"62",x"C1",x"D1",x"58",x"D9",x"E5", -- 0x3BE8
    x"D9",x"CD",x"1F",x"3C",x"E1",x"CD",x"7B",x"3C", -- 0x3BF0
    x"28",x"D6",x"F1",x"32",x"13",x"43",x"C9",x"CD", -- 0x3BF8
    x"1C",x"2B",x"F5",x"CF",x"2C",x"CD",x"1C",x"2B", -- 0x3C00
    x"F5",x"CD",x"7B",x"3C",x"30",x"CA",x"F1",x"32", -- 0x3C08
    x"16",x"43",x"57",x"F1",x"32",x"15",x"43",x"5F", -- 0x3C10
    x"EB",x"D5",x"CD",x"8A",x"3B",x"18",x"D5",x"CD", -- 0x3C18
    x"C6",x"3C",x"DF",x"C8",x"00",x"00",x"D5",x"7B", -- 0x3C20
    x"95",x"DC",x"8B",x"3C",x"CB",x"19",x"CB",x"39", -- 0x3C28
    x"47",x"CB",x"39",x"CB",x"39",x"7A",x"94",x"DC", -- 0x3C30
    x"8B",x"3C",x"CB",x"19",x"37",x"CB",x"19",x"B8", -- 0x3C38
    x"38",x"4D",x"57",x"78",x"5F",x"C5",x"E5",x"7A", -- 0x3C40
    x"4F",x"3E",x"00",x"57",x"47",x"67",x"7B",x"6F", -- 0x3C48
    x"CB",x"25",x"CB",x"14",x"ED",x"42",x"CB",x"21", -- 0x3C50
    x"CB",x"10",x"CB",x"23",x"CB",x"12",x"7C",x"D9", -- 0x3C58
    x"E1",x"C1",x"D1",x"CB",x"27",x"D4",x"A0",x"3C", -- 0x3C60
    x"CD",x"AF",x"3C",x"CD",x"C6",x"3C",x"7A",x"BC", -- 0x3C68
    x"20",x"03",x"7B",x"BD",x"C8",x"D9",x"19",x"7C", -- 0x3C70
    x"D9",x"18",x"E8",x"7E",x"FE",x"BD",x"20",x"0D", -- 0x3C78
    x"23",x"AF",x"C9",x"2B",x"D7",x"3E",x"00",x"C3", -- 0x3C80
    x"4A",x"38",x"00",x"ED",x"44",x"37",x"C9",x"CD", -- 0x3C88
    x"97",x"3C",x"5F",x"78",x"57",x"18",x"AE",x"CB", -- 0x3C90
    x"09",x"CB",x"09",x"CB",x"09",x"CB",x"09",x"C9", -- 0x3C98
    x"CD",x"97",x"3C",x"CD",x"AF",x"3C",x"CD",x"97", -- 0x3CA0
    x"3C",x"D9",x"B7",x"ED",x"42",x"D9",x"C9",x"CB", -- 0x3CA8
    x"79",x"CA",x"BD",x"3C",x"CB",x"71",x"C2",x"BB", -- 0x3CB0
    x"3C",x"24",x"C9",x"25",x"C9",x"CB",x"71",x"C2", -- 0x3CB8
    x"C4",x"3C",x"2C",x"C9",x"2D",x"C9",x"C5",x"D5", -- 0x3CC0
    x"E5",x"7C",x"65",x"6F",x"CD",x"8A",x"3B",x"E1", -- 0x3CC8
    x"D1",x"C1",x"C9",x"11",x"03",x"03",x"18",x"08", -- 0x3CD0
    x"11",x"00",x"00",x"18",x"03",x"11",x"00",x"03", -- 0x3CD8
    x"ED",x"53",x"17",x"43",x"2B",x"D7",x"CD",x"1C", -- 0x3CE0
    x"2B",x"F5",x"CF",x"2C",x"CD",x"1C",x"2B",x"D1", -- 0x3CE8
    x"5F",x"E5",x"C3",x"A2",x"35",x"46",x"23",x"3A", -- 0x3CF0
    x"14",x"43",x"B7",x"28",x"4B",x"4F",x"7E",x"CB", -- 0x3CF8
    x"2F",x"CB",x"2F",x"CB",x"2F",x"CB",x"2F",x"08", -- 0x3D00
    x"3E",x"01",x"08",x"F5",x"CB",x"2F",x"38",x"3D", -- 0x3D08
    x"CB",x"2F",x"38",x"36",x"14",x"C5",x"D5",x"E5", -- 0x3D10
    x"6F",x"3A",x"13",x"43",x"F5",x"7D",x"2A",x"17", -- 0x3D18
    x"43",x"A4",x"AD",x"32",x"13",x"43",x"6A",x"63", -- 0x3D20
    x"CD",x"8A",x"3B",x"F1",x"32",x"13",x"43",x"E1", -- 0x3D28
    x"D1",x"C1",x"F1",x"0D",x"20",x"D5",x"C5",x"08", -- 0x3D30
    x"3D",x"47",x"08",x"04",x"05",x"C1",x"3A",x"14", -- 0x3D38
    x"43",x"4F",x"7E",x"28",x"C6",x"23",x"10",x"AF", -- 0x3D40
    x"E1",x"C9",x"15",x"18",x"C8",x"CB",x"2F",x"38", -- 0x3D48
    x"03",x"1C",x"18",x"C1",x"1D",x"18",x"BE",x"0C", -- 0x3D50
    x"23",x"EB",x"23",x"12",x"13",x"0C",x"C3",x"CC", -- 0x3D58
    x"1B",x"CF",x"28",x"CD",x"C2",x"3F",x"FE",x"03", -- 0x3D60
    x"D2",x"4A",x"1E",x"F5",x"CF",x"2C",x"CD",x"C4", -- 0x3D68
    x"3F",x"FE",x"08",x"30",x"F3",x"3C",x"F5",x"CF", -- 0x3D70
    x"2C",x"CD",x"1C",x"2B",x"B7",x"28",x"3F",x"FE", -- 0x3D78
    x"1E",x"30",x"E5",x"CB",x"27",x"5F",x"16",x"00", -- 0x3D80
    x"CF",x"2C",x"E5",x"21",x"CF",x"3D",x"19",x"5E", -- 0x3D88
    x"23",x"56",x"E1",x"C1",x"05",x"28",x"06",x"CB", -- 0x3D90
    x"3A",x"CB",x"1B",x"10",x"FA",x"F1",x"F5",x"CB", -- 0x3D98
    x"27",x"3C",x"CD",x"2A",x"3E",x"CD",x"1C",x"2B", -- 0x3DA0
    x"FE",x"11",x"30",x"BC",x"D5",x"1E",x"38",x"3E", -- 0x3DA8
    x"07",x"CD",x"32",x"3E",x"D1",x"F1",x"C6",x"08", -- 0x3DB0
    x"CD",x"32",x"3E",x"CF",x"29",x"C9",x"CF",x"2C", -- 0x3DB8
    x"CD",x"1C",x"2B",x"FE",x"11",x"D2",x"4A",x"1E", -- 0x3DC0
    x"F1",x"F1",x"1E",x"00",x"C3",x"B6",x"3D",x"00", -- 0x3DC8
    x"00",x"5D",x"0D",x"E7",x"0B",x"9B",x"0A",x"02", -- 0x3DD0
    x"0A",x"EB",x"08",x"F2",x"07",x"14",x"07",x"9C", -- 0x3DD8
    x"0C",x"3C",x"0B",x"73",x"09",x"6B",x"08",x"80", -- 0x3DE0
    x"07",x"5D",x"0D",x"5D",x"0D",x"5D",x"0D",x"4A", -- 0x3DE8
    x"09",x"90",x"10",x"C0",x"0E",x"24",x"0D",x"68", -- 0x3DF0
    x"0C",x"0C",x"0B",x"D8",x"09",x"C8",x"08",x"A0", -- 0x3DF8
    x"0F",x"EB",x"0D",x"B4",x"0B",x"70",x"0A",x"4A", -- 0x3E00
    x"09",x"48",x"08",x"F6",x"B7",x"C9",x"CB",x"7A", -- 0x3E08
    x"28",x"13",x"CD",x"EF",x"0A",x"7A",x"53",x"1E", -- 0x3E10
    x"00",x"B7",x"1F",x"CB",x"1A",x"CB",x"1B",x"06", -- 0x3E18
    x"91",x"CD",x"69",x"09",x"C9",x"EB",x"CD",x"9A", -- 0x3E20
    x"0A",x"C9",x"47",x"D3",x"F8",x"7A",x"D3",x"F9", -- 0x3E28
    x"05",x"78",x"D3",x"F8",x"7B",x"D3",x"F9",x"C9", -- 0x3E30
    x"AF",x"2B",x"3C",x"08",x"D7",x"CD",x"1C",x"2B", -- 0x3E38
    x"F5",x"2B",x"D7",x"28",x"0C",x"FE",x"2C",x"20", -- 0x3E40
    x"05",x"08",x"FE",x"05",x"38",x"EC",x"C3",x"97", -- 0x3E48
    x"19",x"08",x"FE",x"03",x"38",x"F8",x"3D",x"3D", -- 0x3E50
    x"32",x"1D",x"43",x"11",x"18",x"43",x"47",x"83", -- 0x3E58
    x"5F",x"F1",x"3D",x"FE",x"04",x"D2",x"4A",x"1E", -- 0x3E60
    x"12",x"1B",x"10",x"F5",x"F1",x"FE",x"66",x"30", -- 0x3E68
    x"F4",x"57",x"F1",x"FE",x"A0",x"30",x"EE",x"5F", -- 0x3E70
    x"E5",x"21",x"FF",x"FF",x"E5",x"EB",x"22",x"1E", -- 0x3E78
    x"43",x"CD",x"04",x"3F",x"28",x"06",x"2D",x"3E", -- 0x3E80
    x"FF",x"BD",x"20",x"F5",x"2C",x"7D",x"32",x"20", -- 0x3E88
    x"43",x"2A",x"1E",x"43",x"2C",x"3E",x"A0",x"BD", -- 0x3E90
    x"28",x"05",x"CD",x"04",x"3F",x"20",x"F5",x"2D", -- 0x3E98
    x"7D",x"32",x"21",x"43",x"3A",x"1F",x"43",x"A7", -- 0x3EA0
    x"28",x"0C",x"3D",x"67",x"CD",x"C3",x"3E",x"3A", -- 0x3EA8
    x"1F",x"43",x"FE",x"65",x"28",x"05",x"3C",x"67", -- 0x3EB0
    x"CD",x"C3",x"3E",x"3E",x"FF",x"E1",x"BC",x"20", -- 0x3EB8
    x"BD",x"E1",x"C9",x"0E",x"FF",x"3A",x"20",x"43", -- 0x3EC0
    x"6F",x"3A",x"21",x"43",x"95",x"47",x"04",x"C8", -- 0x3EC8
    x"C5",x"E5",x"CD",x"F1",x"3E",x"E1",x"C1",x"20", -- 0x3ED0
    x"06",x"0E",x"FF",x"2C",x"10",x"F2",x"C9",x"AF", -- 0x3ED8
    x"B9",x"28",x"F8",x"0E",x"02",x"C5",x"CD",x"63", -- 0x3EE0
    x"19",x"C1",x"D1",x"E5",x"D5",x"0E",x"00",x"18", -- 0x3EE8
    x"EA",x"CD",x"3A",x"3F",x"E5",x"21",x"1D",x"43", -- 0x3EF0
    x"46",x"21",x"19",x"43",x"BE",x"28",x"03",x"23", -- 0x3EF8
    x"10",x"FA",x"E1",x"C9",x"E5",x"CD",x"F1",x"3E", -- 0x3F00
    x"F5",x"41",x"3A",x"19",x"43",x"4F",x"C4",x"B0", -- 0x3F08
    x"3B",x"F1",x"E1",x"C9",x"16",x"FE",x"18",x"02", -- 0x3F10
    x"16",x"F7",x"CD",x"87",x"3A",x"6F",x"26",x"00", -- 0x3F18
    x"C9",x"FE",x"91",x"CA",x"F4",x"36",x"FE",x"8A", -- 0x3F20
    x"CA",x"0A",x"37",x"FE",x"80",x"CA",x"61",x"36", -- 0x3F28
    x"C3",x"05",x"25",x"23",x"C3",x"29",x"2C",x"6E", -- 0x3F30
    x"63",x"77",x"7D",x"6C",x"26",x"00",x"54",x"5D", -- 0x3F38
    x"29",x"29",x"19",x"29",x"29",x"29",x"5F",x"CB", -- 0x3F40
    x"3B",x"CB",x"3B",x"16",x"48",x"19",x"E6",x"03", -- 0x3F48
    x"3C",x"4F",x"47",x"7E",x"07",x"07",x"10",x"FC", -- 0x3F50
    x"E6",x"03",x"C9",x"00",x"CF",x"28",x"CD",x"1C", -- 0x3F58
    x"2B",x"F5",x"CF",x"2C",x"CD",x"1C",x"2B",x"F5", -- 0x3F60
    x"CF",x"29",x"D1",x"F1",x"EB",x"D5",x"6F",x"CD", -- 0x3F68
    x"3A",x"3F",x"6F",x"26",x"00",x"CD",x"9A",x"0A", -- 0x3F70
    x"E1",x"C9",x"CA",x"FE",x"27",x"FE",x"FF",x"C2", -- 0x3F78
    x"04",x"25",x"D7",x"23",x"FE",x"82",x"CA",x"0F", -- 0x3F80
    x"3A",x"FE",x"8F",x"28",x"CF",x"FE",x"83",x"CA", -- 0x3F88
    x"1F",x"3A",x"C3",x"21",x"3F",x"CD",x"1C",x"2B", -- 0x3F90
    x"FE",x"10",x"D2",x"4A",x"1E",x"F5",x"CF",x"2C", -- 0x3F98
    x"CD",x"1C",x"2B",x"5F",x"F1",x"C3",x"32",x"3E", -- 0x3FA0
    x"CD",x"C2",x"3F",x"FE",x"04",x"D2",x"4A",x"1E", -- 0x3FA8
    x"E6",x"03",x"07",x"07",x"07",x"47",x"3A",x"1C", -- 0x3FB0
    x"43",x"E6",x"E7",x"B0",x"D3",x"FF",x"32",x"1C", -- 0x3FB8
    x"43",x"C9",x"2B",x"D7",x"CD",x"1C",x"2B",x"3D", -- 0x3FC0
    x"C9",x"CD",x"7A",x"30",x"23",x"CD",x"7A",x"30", -- 0x3FC8
    x"2B",x"C9",x"FE",x"22",x"C2",x"89",x"2B",x"03", -- 0x3FD0
    x"15",x"C8",x"7E",x"FE",x"22",x"23",x"02",x"CA", -- 0x3FD8
    x"89",x"2B",x"18",x"F3",x"2B",x"D7",x"06",x"04", -- 0x3FE0
    x"CA",x"BD",x"38",x"CD",x"C2",x"3F",x"FE",x"04", -- 0x3FE8
    x"D2",x"4A",x"1E",x"E6",x"03",x"0F",x"0F",x"47", -- 0x3FF0
    x"3A",x"1C",x"43",x"E6",x"3F",x"C3",x"C2",x"38"  -- 0x3FF8
  );

begin

  p_rom : process
  begin
    wait until rising_edge(CLK);
     DATA <= ROM(to_integer(unsigned(ADDR)));
  end process;
end RTL;
